PK   ��W�� ��0  ��    cirkitFile.json�}o�F��ߊ����v��O���lr �3��$�������<\~y�.J�%Q���oM��������b����.�v�,jog�b��~j������J�.(��������n~;[-f�/˻._����V�޵Q�l˦Z�}f���2��(��.rq�DyW&Q�Q^'&�e����\������H�`f$f�*�Y,f�*��3H�̉�
f���
f���
f���
f���
fV��
>F��X�S B�<V�<X�%<�<\�%<�<`�%<�<d�%<�<h�%<�<l�%<�<p�%<�<t�%��J;��B;��0Д��X;��B;��B;��B;��B;��B;��B;�>'��N�����N�����N��� ����i�S,�)�S,�)�S,�)�S,�)�S,�)�S,afN;��B;��B;��B;��0�)��N;��B;��B;��B;��B;�f��c�X�S�c�X�S�c�X�S�c�X�S�c�X�S �cg"��b	O!��b	O!��b	O!��b	3K�S,�)�S,�)�s q���]F�r~����nqS.�_���H���{�a�Kg� �v��݀�I�^�x��moW3�Uy�*U�Ƒ��:*�:J��RV�6��%�a�k�kv(a���bmg����ѐ��w��>s���a��#,��`m�`m7�;�c�5i�u�Ig�VZFE֘�x+).����{b~x�5{�5;���tf�am�am�#,���X��X�A�Kgf�v�vP:���k���<8����_���A��ǯ����k�|��^���6X>���`���,�;6r�]S��+"Sق��8*����͋�(�iәf�Nq��`���oW��NV�|������',X>���`���,���]|�������|�� <#N]�|���`��S,��x��~�G2�g2��%�.18u����Wˀ�N]�|t�O�v�	m�ebp.��#0�v���`�������2X>��
3�������|f/�B��e�|��C�9d_d�y��EX>���F���y���|�*l?p^��#0�'����}5p^d�y��EX>��^�������|��l?p.��#0�����`���+����2X>��Zu�������|��k?�?�|��� `���,�����~���G`>�� �8������I��^��^��?8�p���G`>���8�����k����?�|��)`���,�����~���G`>�T��_�?�|��;`���,���:�~���GG��Ԟ��E[k˨,�*ru�GU�tQ�Y��:IM>3�G�	8uI�����|\�	l?p�2�;�jA�WR�s�z����%�Aw�x�?8aJ�	SN��|�Lߴ�I�6�j�ȵTEE�Ū��LKm��N\�{j\�lzp���#0WY��ka��������ZX>�qe;��Rp���#0����ka�������ZX>:�����(lb�&3r��VmE�����#gr?4q����X��e~0�xd��H���ERU&o��U}�a���]�6uѕ]��<���?��P�Kٻ���� A��IR='�},�NF�3Ӻ��ʨ�s�%gI�NM��4+���J�,�?+O�������k�N.�Uv��?���4����t�Dtl+:�(��(6Ģn����c�����a�NG����m��a��ݭlw'�P+���A�qX�~���pXq0�+@�q�v�q�v�q�n�$���ݝ���n|�v��B?|_v��B�|�u���d&~�
�cI`С��:�#%A�a�{l�:b�{l�:R�{l�:B�{l�:2�{l�:J�[]����;���Xv��49%:����S�?ѧ��t��O�ey�.	|sC8<����r�1��O��]����y�$d@8�*	��#������	�<6&��y�w
�$7Z.94	��B�=�d<
�Ċ�DlH��r%Ws,v��"�]i��B����dgr�|���=�l��Ջ�����oO��?���忙�����O���_zHȰ`�@B��
C2<�!	�����ϐb�@B�'J1D !�s�"����\H��3Ġ��ڸ����(%�ώ��`��`��d�Y|,~,���L������(%�?1��x��(%�?G1��߸8,�ǰ8�R2��,�ǰ8�R2��,�ǰ8�R2��",�ǰ8�R2��%P:���QJ\�Ƅ�I�M��⸅�q���1�⸅�q����1�⸅�q��@�1�⸃�q���1�⸃�q����1���q��8�`q����`L�8�`q��e�`L�8�`q���`�~`q<��q���1��x��(%�Yc�=��=ބ���QJ\����	,����L�	�SXG)q9,���8>�4�l�a��j_� �J*���j_Sī�:d��s�*Ю�U9�@�j��
���7����:x׫R^|���Y��!Ʈ�1�`%VsX��
��_5X�EŮ��1v�`%V3;�FW�U��TX��J!\hWVRa5���pU�]5XI���	�It2.Zҡ�w�ul��uiВ-���c[��K��th�]s��d_*��Ck�j6!m�����W�r[�I�H'S�%Z^àc[�LL��thy-��mu�1Zҡ�5%:����ThI������V'+S�%Z^��`A'/S�%Z^��c[��L��thy͕�m���)=���b��,���ThI������V'/S��c���,���b��L��thyM��mu�2Zҡ嵕:����ThI��׈��V'/S�%Z^�c[��L����"�2���Y��L��thy�mu�2Zҡ�5�:����ThI��ׂ��V�mE��u�2���Y��L��thym��mu�2Zҡ�:����ThI��k%��V'/S�%Z���c[��L��th�v��mu�2Zҡ�*�u:y�
-��r-���e*��C�5Qtl����В-�vѱ�N^�BK:�\�FǶJ+ɔ����eN'/s:y�
-��r� ���e*��C˵�tl����В-�pұ�N^�BK:�\�JǶ:y�
-��rM-�&:y�
-��rm0���e*��Ck��"���N^�B;��&�z���%:y�
-��r�9���eGh!�(�j|(�P��T�C'/;��,ҶCZ�mu�D'/Kt�2Zҡ嚌:����ThI��kK��V'/S�%Z���b�T'/S�%Z���c[��L��th��g������Th��v>��M�f�W�:�@��M�涱�@%���=>,��� ,}��+�
T6խ�*#��'��T���2R�y�׍�i�*���ܺ�$�̦r��B"��o�cK��[�؅�$���*%Nr�?`�u�f�er�ԩ��T��\��Q��Udl^4EQgM��}4~��H!�*#��'�X���`�2R��Jz.���VA*g�U���`�u ��x�����`�w�;�Se0<���2���T���1i&�z����t+a2g��0��\�&c���a2�\�&��G��`�ܱ��N��8-�8Æ��^\Pc�D#�����O���IU�[%�]�˘(/r�M]te׺<�֣��=f�
��E[k˨,�ʫtyTIUq����Ij�5�X��� ��\�
R9�V�j+*MԵU9�{=�Qj(��5Y^n�r*�R�s�v�Cb�ue��y�Ϩ�3rM��iQ�iV4�]��J*�T�\R�*/\e��ژ�����)�������jm��ˉ�:H��]� ��C� {�h�ʤi�D��6u-UQQ�IT�MgZj۴�L���SA*g��r�.A*�v�������U�j/_��$;�{Dl���a�,ov���$dz�C�@B���"����B2}!	�>����L��C�@B���!D !��@�@B�������z6"qQ�aq�`��d֓6&X�&X�F)��t�	�	�QJf=хa��p�q��YO�a�`q<��q��YOb�p�o� �cXG)��(�	�cXG)���,�	�cXG)���1�	�cXG)���6&��q��(%.\c�ͤ�R`q���8J����`q���8J�Z��`q���8J�(��`q���8J����`q���8J����ps�IqXw�8�R�B0&Xw�8�R��0&Xw�8�R�B�G?�8���8J��Ø`q<��q�/Ć1�n�o��x��(%^0c����QJ�@���),���xA �	�SXS���o�x��^�P%VRa5���Q�*Ю���jf�E�hU�]5XI����|Ъ@�j��
�ϻT�:����+���q��]�{ �`%V?FQ��v����jf��=hU�]5XI���E{Ъ@�j��
��
��U�v�`%V~'X'1�ɸThI���mֱ�R֥�v��]��x�N�BK:�����mu�/Zҡ�w�ul����В-���c[�,L��thy��mu21Zҡ�:����ThI��ה��V'#S�%Z^�c[��L��thy��΃��L��thy���mu�2Zҡ�5W:�Uz"��HL'/�u�X'/S�%Z^�c[��L��thy-��mu�2Zҡ�5�:����ThI���V��V'/S�%Z^#�c[��L��thy���mu�2Zҡ�5�:/&��e*��C�k�ul����В-��ֱ�N^�BK:��\ǶJo+*�����Y�����e*��C�k�ul����В-�б�N^�BK:�\+AǶ:y�
-��r����e*��C˵+tl����В-��P�����ThI��k���V'/S�%Z���c[��L��th����mu�2Zҡ�5:�UZI���L'/s:y����ThI��k��V'/S�%Z�}�c[��L��th����mu�2Zҡ�ZT:����ThI��kj��6���ThI��k���V'/S�%Z�q�c[��L��th�V��mu�2Zҡ�s:����ThI��k���V�ʇR���,�����L��th����mu�2Zҡ嚌:����ThI��kK��V'/S�%Z���b�T'/S�%Z���c[��L��th�f��mu�2Z
�}�T�mM�gEq����Q�5&2iݕ�	Un�;�UFj�NT�&;Qe���D����UFjeOT�n=Qe��D��
�UFj>O�:��b�w죯Se0�;�iթ2���L�:5]�����8*����͋�(�i���*H���R9{��T�^� ���:H��R�\��*H�l�
R9�¼��=��d0�{>X��`<��>�<U��c�!��0^<��ߩ2/���T��}�v�Ƌ�>;U��ca���b�x�S�;2ERU&o��U����"wQ��EWv���,`T�r��,��Z[Fe�T^�ˣ�H���K6�NR��g	R������T��ە�ڊJumUG��^��u��jcM��v	R9k�̴.�2j��gT��&J��4+Ӟg	R9��*/\e��ژ�����)�������jmr�%H�r�_�T��K�V&M�$����k����L��l:�Rۦm��J��Y����K�ʮ]~���e5�7��l��r���˟���~vwS�m3���˦]^���[A�x�]=��$%Im�O�GP�9����iрSb�8=~����yKn?�����d��{�ءCz�y��<t�l�؁]�h|<r���\4������I�R\�u2���{(�����H����<|�&髍�y�PG�2�	r��1����$0W�<�yd��8��:��PE�ڣ�f`f�p�g����b���#��5I�K�����HF��֟n��s���m�e���'����ͱ��[���e����"i/'@��'���t�$�����F'� +Hs|���>�
Ҍ`i����'	��4@O����?�<!������@�N!��MR�/#z�B>,AOY�o6�̅<�q�}�c����]B�)H�?�����I��.�}����Nxnh�>fy� ��p<}��4�{���'	� 9�p"l�g��P�l淋���\��/��躵�l��=̛��=�Z�~���mC�[�k1�]ܩ$�0�k5B
���_�R�%L�Z��B,a�B
���@)��_@!�K�~��B,a�B
����)�f��D��>� T�a�k`��J� *�0�U8R@%@ �k��: ) � ��5�z%��Oc@<�k��Z()b<���i��r�^�%� ��O�f��L���1 ��5�zI��Oc@<�k���:i*	��O���< "�G���xj�T���)p ��S��
���O��]%  �:@<�k��z �x� �T��߁p �L���x� �T���� p ��S�����O��� ��> �&�x*���� @<M �T������P��P�x� �\��M8 �4�S��1p �i
��r��� ��O��k�j&���EgEz�#0�9|���߀����&1�2NbN,���l���~X������e�?��М�O�O�G`>s��$Rb�߾���5,X\?h �s�%�9�|�3��Gcpz�a��gf���� ��������A��#0�Ԉm��0!�	��L��)��Є�2)چ�<LHhB~mCt�&$4��[#��!:A��2>ъ/~mRt�&$4!�K��!:Q���G����		M�ﰣm�NX���&����6D'-`BB����6:m���=�m�N[���&�5h������Ӗ����LHhB�W�	cCt�&֝�-�'��mRt�&$4!/YB����		M�˭�6D�-`BB�R1��i��Єf�4Ɔ�L8�F��b,:���,LHhB^m��!:���WJ�m��b���&�U�h�_��)��b,:���,LHhB^]��!:m��W�m�N[���&�U�h��0!�	yE6چ�LHhB^M��!:m��Wm��y
��Є��mCt�&$4!W @����		M���6D�)`BBr���X��X�y�C�)���		M�7�6D�)`BBr���y
��Є\�mCt�&$4!WiA����		M�f�6L�y
��Є\mCt�&$4���BƆ�<L8�(��Q��˧\�mRt�&$4�|=*���pߋ���C���������g���1):�I�I͐� �IM��qt���s0!�	��چ�LHhB����!:������m��s0!�	�bچ�LHhB��]d��9�p�)�A����O�<�T�쓿9�w2��Ɏ|�2�����BM��'�.�I�;��
�ܠ����P'�?�\:�3%G�
}�H����mR��лM&����%zC�6������H����������%`'�o���G� �A%������+h��+h��+̻��)���73�
H=t��ʩR�~r����_b�*Po��aFX�� ��2L/���;�͎t;azG�ّn1L�H7;�m���fG�az�nv�	�����9��� �1���T�S��H���m���0Q^�.j���ʮuy�������960(�,�֖QY6����*�.��ҟ�����G�h�?�䎄�o�;-F�!H�H�ɇ+[��&�ڪ��ɽ���(5��ƚ,/��n,��;����.3�K����:o�ɖ|����<-�8͊ƴ��Fl$w��F�몼p��*kcv�:*�:�	��'���ߍ�l�����$wbp����h�Wj�ʤi�D��w-UQQ�IT�MgZj۴=6-4��k�o��N+h�#�J.��|��7��b���/_�v��^����M�>���!��.����9�����콯7CN�E��T���|ۀ�zL�_ܾw��F�o�> �A&�=��$�=b�#�=b�#�=,��/��Y���!�tx�~ǐH�w��೷C�x-����=�a퀷��o�y9s��w}~?'J!�4$�����XB#}���Շ!������2�s#t�����o��H��fT�#8��:��·�!N&��h����E����p
�u$O���Ţ��8$�C���8�e�C���8���Y5��؁O1%�%3���_d����C���2ӏpX�O�{Xqi�;��� �tc�R����!�X�g��ܝ=�cf�"8{�rc�W�����L<�{�I^�u^��^�f�0c}W����u�!�h�.M}��6��N�jY�nʪ��d���|q�u��`3l��&n�7���&��d���f�nJ6���t�)n�6���|�)n*6���&�Z���Gs�A[{�� �5-B[���$�5	mB[���(�5
�B[���,�5�o��o��?���.����_���77����o���f~���wB�������C;��q����Sx��g���x����\�^����o���v������w��?|o{3ܯ��[�ݖ?�y���O����o�_��s��۹�����a���O��勮��o���v������i[���0_��動��f���}��z��l�� v��|�zQ-V ��#�|5_x;|�I�k�P�o�ޜ镵�:q�Q��OoZ�}�%.��.�,���,#�Q��3��[�f~��v�����Uy[��	����\,��ڕk������|����i7�y���0Y��k��*&s�
���4{w��ׅ�&M�?�цy|��>-ˊ���\g'�h������Dv���Y��H{#6lt�\\$���.)����ɒ������~�"K���oG��y�ܸGB��/iBG�%T<�I�����X�K�k[����ǵ.����?�Wd#]l�a���ohɦ��Y+.6���vi/�����ekB�6g��5,ւ�6����~�ӟJj�3�������WoV�|�vy��k�����]il���������y��.౉2��v"}v�\v���e�nl�mS%��(K��,s��Qk���dI�o������065��o�������nǁ���������v��x�w��{�������{jmwD�~}�1����	��'������m�G�1c�P1�e�������}��>4�ρu���ʲ�V顖;ڬ�Z�6���l>���*����oX�!^u���]^��]sw���������.����7�/y[�[&)��Tf��1EU��KlV��Z?r�۷���,|T�b��������w��m�1B�SȪ�c�̸�K��ŵ������g�i�<K"��W~���Q��;�+�.����=�����a�{P�2�2�#��{ꪳY��mڦ&��,]������-K|�m��6 =�ɧ?�o��&!�V��*��8�6y�[:i�tuc]M]�g�O��r�zu���\�WT�Yd�ƫXj��*�(ɛ��|�^t�����ݥi}Gn��FMGq����As���)�IW�y���y~��]y۴��9���	�?��궗��n�z���~���_�6�f�\}�4���~#���'���7�׺�{�Wn��(��t�_����Ⱥ�Q�fIY%qV�z̽�(.��4J��[2��|n�5ISdq��Q����;ʛ�n:���6�M�|�o��u�R5�^6�\Wm�I������f7u.�����{��~w�oM��oۋ��go>��ͫ׳�/�����w���}���o/�Φ���웗_��x���>�����]��^��o��쳿�t��ly�ɛ���g��_�������x��������j��������_)��oW��|'����6�����6��?3�%�)=�%�[����l�G�d��f��F-?��Ŋ���?-���}�z���C����..�~��k�o���_.>�18��x��.>��l�х?�7>3�x`��ֿ^��Y����]��M����C;\]����o���Ï���[$�Q<���N#��L�f�h{�������C�}7�m��l�#D[����_�j{��Յ���s�o��k��j/_�io���8�_�f��|U޼n����6,[�
ۓ��	�{Η|O���f�7{����Z�����^|���˱���>�w_�׾%�����b�_�s����և���<��{�gS�}Xޮ�B8�)[0�8�	[<°,�0�a}t�P�������9�O..Jvq�Vܩ�����m����8�V����.���	..�����?�}���}��Qv�wo�]��.��]�6W{���m�F�^������e��[����j���?:��������W; �5	`G���SaNt�0�f޿g�|���������O�����>8�4?�����-���n=P�����}�Q�30����~�Z��Ay���N��~b�o����g%~x��o��u�"�%sz��q�67߱6�~&���w�2���=���G3_O�p/����/ϡ^��"~e���^<���#��	�#�7�M[���j=�f�.�)�������f�y�gT���r�ܕK��$.2c����\�>aH�N��6e�|��.^�6�O{������'�\�.�v�l��gv��3�6�l�&�Q��e�S�����$��\V�C�?�2|�>���i�,>x��s8�Mē81O��O(�QmDI�'ysW.����-�3Rg��Sg7����+����d;���T��dEm�dQCu�e�:�ʬ��m���=����ꁃd�Lp�?������zOp�)�v�+k
�=�<��l_�O��̇�M���e���VM��2�?��8��i�\��u�&��<u,��YT�-L�6Q��>�4޹��-��Ω횮��:����#AȱK���J����ss��L���%�#�������=o�:KТ����%�S��d�X�,��7Jn�ỉm��JWQ�]�-��+
��5J�f���&��x�_F����L�vY^��1i�%haT�Q2{�p��ߎkmqM����֟C~탯�����d?l�&��%W���&K��o�l/�]gy����_�4!��C67�6�*��565q�H���,��}�W$�iͣi=*]�4N���[tc�m�F�nL�y�!�t�k�^���:�C�< ��L�����d�o���;�����5���ߨH�w@8�<oV?��i*�����?���o�����k2I�*��ο��Wy�>ek>y|�����~�Ǽ���>����T��#���r�����,Y�����\�$t�$��+��dn��Za+�z�e��(���w��Y�7��^�'��]�k��oxÛ�/��__|���?�~�������H��m����V�C��V�c��x�w>���{ݾ��ҁb�s ;І�@�,�w�;�~+\#��~���@'[w��?��@ak\O��x�k�CM`�'�D{Jב`/|�����k�wֈl|��w�V c}�=�w&�"}�����9PZ���V�4;�>��K
����A]R�B�p7��'M�x�w�y��W~��ݝkJ�!�]��\:�հ�<�H��C�T|����Hg�������������K��4��(Ѝ�I:[@�(�Q�v��F	&=�8���F"M6�Q��h̖P7:5R�\o�Fg��������n�n�C��;kީ��}h�X��F�F�F�F{�N�Q`��q���Y�#����:Rt�	s�S�`�������hoډ�Q`�1�4�Up�F��+�b�tXm"�b����s�ASл�����PƜiu���e�u�%+�y�%�����&���C�"w|".yF��h`C�0�Yc�I�~aU���~�3��&�"����N�3�}�={z�w����'���9����a��Cy��'�Ö�ZdP�9(/�}Ό�1�S{#4g��*�3�3� ^V��!�SklJ���z[	#__��2'2��v��xQX��G�/'
���zv��Y�p:�=Ue9p��ؽ���F������6�yW{�����ٟ�ۦ����m�Լ� ��m�B�D\�:�9(Uz΅0����1��Nv�T+h��y��C���z�A9Xp����3^�yz}w��©9���*�|g��;a�y�I�s}g+2����n�����Z�.�w�� 6a���I�3�k&�"sn�t�����������*{�O��
+k��̐3�7Gh�1���[=�49�&pX+�ǡ3�ƞN�]��!�nxPvV����5�n����i����ː�\σvI�{}G���fO��N'�IW6�Dس밂�`�~r=�nz^�X�69���kZx���{�5s��Ĺ���Kc�AzQ�c̰/��(�)��g�mm��;��5��^��0*���yx��Ɔ���n	cG����;���O_��viд� �	� 6�}f
3���S��t�^��ӱ��h�凃Lf����?S�I�~��Ytj�ｴ��phd����Р���x�����U�U�j������;�}������W��Cy���Ǘ��G�����/��PK   ��W`�����  (�  /   images/a675022d-8297-46f2-a9f0-ef789ec00656.png�ZSs%�<'9�������ƶ�ll�X'۶m��ƶ��݇�'�T�K��tMW�TM���"<.<  @��U  ��X��t.T  � �"���������/j�(n� nADB��O@�_NȀ��Q��5��!5��)!����1�������-����sRJ$	D�ׯ/tL8^DQK����z���ӽ����Wd1S<¯�wFfvNhV9DY;x!cXvuh&)����OD6%,l<N%>���Wa^U4zћۛ�����d(
�ǧGV6Vtfi�,��H<W�4�ș��Y�ܗ���<|}a(�K���w���R�c����f:8�}yy��ҽ��¤�^]]�64���XX�%tY����b�����FP=:��&�$&!�ϧ�����ю.��EF��������xb����R���)�3���������?x���յupy%��o-m��=�a��p���u	]�[��u;pl�M�-p��-��c{{���呌{�C�I8q�����<y���.V�;�%mSXR��+K�)���G�S�����K��_����b���>���C�ޔ�؍����Ƿ������ёOR���CHQ�]N��g��oQ�҉HB}��{zixySB�R������IBy���52��ɳ}~���od�
1��9�c��7J��o��rl���ӇsPDXjN�꾴�~ra�`���W��\Hv���������"��Ĭ�֫'8.y��A�,���5>�XÅJF�5v��+P�1�KÄ!|�,0qn笭op~gg��bf���k����#�M�Զ[J�@�^��id[�0�N���o�<�B(�S�wA=P�*�n��"!�m^$�#�7@�?�8+P��)  H�
������Y�;��B�`�"@X^���U��"Oa��7W�*�S��BL�>��6gaLV���GJ���������zm=wD�{�J|\T択�Fob�P�t�ɨ V��b���h[�Qבץ�t�M-��e���?:x�o4A�/z�$�JTF�TY5�@<>H�Y�j�	�څ�q�����:fqՏ������y�~>\`�������ԗ�Z�&�\�i�r�n��\���X�h���uԮ37�c��LΔN�m3��v<����Z��X��r�%��|<��c{g�k�mc�T�B�"��a#�`z�J�sD}�$�G{��IC-ص\jF����r)�f��0��\vg�d_�!hJ�O�r��1� �`P�sCX0�̴	�Zt4���(�l#z�wm��`;m���x?
�X�S���%W����O�*P(@�51��nh)BF�*5:���@#�LZ��Q�Q�B��ʢx���Ew Y��\��A���8m���a���f���'���m$�J� N�)��� -&-t�������ȡz�Q�!*/Vs�m�Z�-�n^I��#�����j��>u}��T��%z]��}�x�E���4�ZJ4ŗ��v=��$�E�r)o��]%7cRC����Z�j��:?v,�I�����]�Հ�9�2=�����L�2�����A�3��xrm�J�i�����7XxS���k��bD�d:�:�&t�8���>�p�N�Rs�bg��^\Џ�����yP�Ym��H�52�F�󼺽�չ��ڴ&̐ޘ,��Q..�W�,��|{���5R��B���w��@���䯮O��{dzQ����j�F�p�4����)mA�9|~��˙p/�.�K�6�Vy�[��,�+�bn��W��P6�j�O�uqT�Pm��7����Х�F��Q"廾����v>b�D)��ܭO#K��Ȳz��>_qo���7�[��~�N����/�c��,�+��?=���׶LY�����?5����?�*��I|Jk`��{I��p��<��C��:��rĪ�G�!*+t&-B.-��פ��ѕg܇iJ|�]����s%��|�;�d�~uU"���~�U��m�1zs�D�A�������������l6�+�~�9�����}ou�4���~F��kX�r��~t���i�^�,���'Q���C%sֈ����^�HC��-���Z����u�̽}I#������~I%^�"��`|\H�|����*..�����a��K��wѬb��.ƎY3��q[Nq2)>��S7eִKߟe��D/˼@�<J��3��=GN�SP��f��d�I���U�֎C�����u�G�'����x��Kۛ��	=��.��'���3������Gb��N?c뭞�TY[ʄԪ̬��|][>������F}ׂv�[I�O���2�F��"xUuu�#	���Nf�e6.B8���%���/�t�u�}�/���q,%R�6�����hx|��U���666�F��닪H�W�6�x]^?��TY��q���������.r綶|�ۼ��ۻ�|?w&�7�\Ύ�e����(�M���6,X�}�W8
-�[U�iR�X��~W�'�DW��^<kn�V��1D��"��������E.�;W���7��ND������6��%�1�7,%���*�Èc��}�po��:5{㌿�g�b�7�{&�Ӎ�]3\�'G���~G�o!gd�����F������Le��<�.B���ă��
&�N#K��_�M��	D�����:.�-�lD�<l���"��@��/���k�a��'ZNnH���"�&�pz��e���g��hCl�{�BQ�l��P����t=�>}t��\�Y6�u���a�:������u�kC��nx��:�"?47�>��\Wlw���1��0�����B����3&'MӖ/ci�W��7�4�yW&�)���xt�0�A2!v-�IÊ�ul�d�P9���h��bt�p7f��.fim���`E���z��w�[w�����ǟ}�`�\��4�@�oep�d�j"���f����}�}[.�?��v0��>�Zu��K��K�������x.d���d�|#""r+��z�oi)�NqgM�@��XQ��J(w�vhkk��m�L��D�.@�D�E��:�?t������+�j�Wυ�Ǆ���7�h�'����`S�e�)[����꯿ {L�u�ϙ���b(��N��U"y��O:��k�	�G���-�9-pן��,&���=ŝ��5�1`�ߥ��3xϷuu�-x�����N�����,���������C�I3����$`��]/��n��+��V�εo8���L��ʯp��9aʣ���+�8��9::���{OO�L����A��}یc0H��A����DLO���Z���4'Jo�ʩE�g�':�6���v�.�.��W���)I`��N��c�������9V��ӆ��6�LcC��v<*�y2~	�c�&�+�y5`�K�)E$��C<�V�4�����۳R��]���	|���9SDp<=y��r�.	ō��Tx� b.���)+.�ٴQ���ȸ9U���	 3���J�����a��B�I��w0cB�(�-;-m��vz��1��S}"���n3�3��#�sY�:W=�U������ �8�J٘���M;��,Q�GC��I�~�Qfu`�D�0vwv�����bc�_�s��:3�	�+T��I��~q!��P�@��n|Ęi:_X7��2%~�O�TaU/(5� W�^�>�C����)R3����7x��F吏"��e��xe�ǽ��	0��Ǹ����t�CF9�Å��nC_�}���W��Oe�y�ܭa}�\{ ���2j�����^��(���Ʈjj!�l�-D��M��A����j=؈���Pj�#%�J�Xk���"f[##�R���I9:;9!Ae`3�� ��#��ezF������!��$; W�ԛ��3�5	�M�����6+#!�\����#��l��L:���+(�y´�;#�,u�g�������%�!DY2���Ts;�3�X�Q���k����OC%���LG���n1�;7<���c��U�����,V���k��N�B̏$��wn�_���;���˥6qn�u{�y��j����YS)�O�$Ts��ұ�I����wzFJWy���O����8
y�%��/�E�;�~��� ��/>,�ǂ2����JI7%{�9!���׸|�@���ڂ9�7Jb���倣��LLL/X��mZz ito�HACP�~X�8��$#�h��/JT��w�\�m��<J|��[�Zk�^%~������u�|8�I����[��t�&�2	��H&{��:�$h�J�R�f�7xYtWշ�خ�W�T��;�.��`.�_J �<(�X����"䭯��~��n��v�i[�����Z��3_��8)��]��G4��#/��YK�=������f�~}s�yPT�Ѫf����+9d�$���C��spO��}�ނG(rDh�	f����V6ݏ�|gL)6;p�RA*;۷*�h�#\��IT�l8X��>�������m���T!�}o�K��F��7�,����!݆�ڮ���tt�C��"�t�:��Zr�M6�U{���R\	��{����v�8M�
�����`���Hw�WL�n�����<<���C]4����n(<�}[#������
3E-�oB�ڂ��	\�o9�\�s9�.z?0P����GYY�mLi��4�m�J%̏*�$g��f��S�Ӆ�Q�6���W}t�&!~���g��r�1s����B��^�E������ײ`q��4�^+�K�]���.�=<Z |��|���L�58��_g�ma�g�M 	�6�aV�ňD�A�K&�65YG�>��7������?��3����'׃�'M��~�|��ޏ?�E,�����J����(z����A��D�Ё�Ԋ� ��)�B/нp(\��"������l�O���`��܀��:?al"�`.ؽ���,4��B�)C��O@:"'��Ot�N�|]�?Qk����j��el^^^`��Z#����Gx�u9���=]��ο�L&�c�fKm��A\�;�*�pph�F9���^��)\@ҔUo�l'�(��*/=!�4F�/M�f{�M8%�F�GAe�J�J�"���q�Y�����rk*��;z������d�1b�����7��
��mļ��ɝ�-�D�v��>�/z�9�op�{I����NR��{��_"��C�I��5=�a����R��rM��}<�L�8K`YC`�l�r�1�)gdrls�ZRA�C��*��a�7م�� �S=B�2[?��kw�Tm�8:΁�g�������u�PnD9X\\8}��v�'�O�vDoL�D�Z<�Q?'c �����E�;����pEa�:*�K.� F"(���k�濁:!a�����)�<&f���t���"��w��-�K�
[�
���k�9ض\!R����J<��~��B�����v�ϸ6��<��%��i9z�����'[�	�+��J>��wv��f#f� b��U�z����5�VDi�,Hb t�x�
��y��b�b� n)R��R�l㫁M�D#?l�#nJ I���(��b�mAc����u;�[E�w��o�cEz!u��da�1�c�{^?13mx?ʟ�Cv��j�O�X���dY��xC4���ئ��7q�\?��e��������53Q��D�\[ȍ�Mb���a
n��68��$�j��ׇ����
u�{�����˒4NG]���fzq����k`�gܿ��ﯔj�IYs|GJv�V�y�^��A;:��f�++;C�d�&�ʰE�����9h�si����(����僳�q�+Q��P+q�� �U_��U����H�+	��}!eOE:���i
�CECC���G�4���0rc.�D�C&�5�˃a�=�����F<@��g6��&�!*��<�|xx��399آ�dץAC����Ȥ�;�u�J�cy�c5��WiҢ��L�ӷ�]����y�@�CU�w������)KKW��+梇��X��Y�Q�-��5N�%� �2�ɛ!L�F���Pv�[?��v˚�@3��dZ���GǓ2[M1_�*���������a��`|�d�����mP�R�,����/�y�q(�ȣ�T��y�g�i�~6ܽ]d���j~�a����"��Q�-�i�u#�j:ԧ1l�>�!	J��  n�$���P
,�8B�_�VEs��+l�&�C��S������p���&�RKT���z*��M|�s�^�%���tuO|n^��F�!t�f�J60O#��ьO�<�Mu��Iz��;j��,�lV��L�l��u�h{:'.�"ih�@�y�NWzRȱ���| ��!�� p]���L݉������� *�+�^����UU	p��Չ��=�D���ny���S_��e�n��o	¿�U-��*�'Cc��d��[�&&i��ֹ��v�T�톣v/����t��P����S�It����� _��B��Z��R;�*lBLi;N�(������Y�BY0Z��F-6f>i�|�"� b��er��m����d�oO۞�2[�l�(*A��0qD�m��2�\^ƞ>�T�ʨ�(y�w�/ �7*�S�2Y��j��nG�ҽw%�ʬ�M(����� ƺ�p/�^��C��S����A��K_��J�(\�/U�>�0*� ���e�R,�GLCu(25�'�mO@���V���$`�}���(񨔙:J���J	M_��D�C>?�m���-�P9a}���̩�)�ѣ�퓼%��p�"-|E��ϱ�pQ1Ĉ��)j��1��|A`��98��JӺ����,=��r��\��k���~�x�hhpvwx�z �|W,��*�bױ�u��Vy�w ���KSKMM�_M�&0�=;�@������̏���*x�3x�m��|	)r�Q+��F%�ޫ-��ۃ?p���uŃ��А��Z8)���P��k�vʨ������i�ٞP��S�5L{��GG�Z���V��*)cv�a��?.��!ɽ��-��� �J�"W��\ GȊ�J̀��RV����L�rW6�2�������g��#�M�?�E�� �`�/̞f��o�V�מ�O9�2��n�ff�� ����G��lm/�Ի�R��~:��!���d�]�ITM�+W��3����n;82�)v��l���!i�y�}�m�_�n���0Nq÷��gxy�˷�"=��{�x��H��Y���@�?%S���w�����"�'��
�kpϒ�H5�:�����
!E���T�e�(G�W4�Z��a�z.M��"7�I�����-	�P����3k�Y�>:��@��}�/��Upj�A��%$	-��Ţ6)(;!� ����ԜH��H⺓"`4W��_Hp�D���9ǐ��$�_��˛g�j����(x�L���8߀Q��~��y{��Ч��nW�cG����| !�"/sEP.fw��L���s�۞|��f������$ \c�{����-g��n/��)��q����4�� ���}||�Xz�9x�.d��x�N�W�U�C��b��&���=&�+�����f�6�%��9���nb4
���(�4���by��D�a�y�YK��~/�Y��&<ڙ�Q�7�Ο���s����x<w}�~�3`B�� ���W[���'4�&a4�!*a�TK:S8��Cin�1�lJN�M�������qb>�~�z���m�c�������Λe�'u���c.~4�����_�s\xqe��e=1EX�:���
�A��0K�=)^D1��b%j�r�h~��[��c���S)C����*>ɮ�;��/�n�8^�O�3G�tA/�J-��LN¤O�_�͈�233�ٷ����XK�^����`��b_��E�]t:��Ą��D#���<ۛR�3ǡp�sgKn"6 w�
֡@1�#QY�O7!��::��
Qع����b�L�U]��)�(�Pk�X5hFV�p�YX?w{+?G�*-]����(^Qa�[4�>j�{o��&��֔:�)��2�.3�ݒ������7���ě5g
M
}r*���'j�e[�ՠ�����=OD_ ��C���j�)�������U��-��Y�[��X ���/!g�*���6�hy�Q��߻��~�H<wF�ڨI����v���u�[��nq?@0v����w/�.�'�`�,t��9=i��D Ir��E����WpLr&��K��G��8w#���/>���܂�g������
������;j�$ɑ�Q�C>>a����絬ы��B��T���!��%�����Շ���� "1I�׀�xso&6�u�]go�B	��2�6UPJ">_��6u&DtN��\���o���_�o|#�K���d�+�#�尧�H�jUg�H�4s�襷q�����x��!�:y��~��|�ob�|Hz�8���
K�Bh�=�SM"���H�P��II?5���O/y��&�/��})?i��"�h���Wy�,��3��%��n����0��'/��l��7N$�-�w�ݬ,A�Iʟ20qcd�w&V���ܷ �;Q�/��[I�����N��(;f��@<��#�f��Ry�>M ����8%�������������&7���# 1��|n�42|;����u˞��qf��7ZE��vN��d⑫A��L������^�X����ژ��	[1�p��N��h<�_��yG��*�Ia��y^�$km'�*� Lg*K�0��n��
>F/	>�:��� 7._�,X	�HR�����)��t!�kQ�Bz��%͸^J֓�S������;��X�����P~�]���ǺQ='v	��ۓ��?�P��ZLrۛ�%#@�D�
��GR���CՅT��@�f!���5ۈ�����MGS4վ���/��ZYMqfrC_OUiK	>c�ց)Qz'1cJ���;��܈�CpƞǑ!.�7�9�սI�q����xŘ���R+�]_�gQX�ފ)Tb�l���� �l��r�l��{��Ex���!�v� ��#�����n5�SpvG�Ce����V�k��Q��~��u��i���_��H�����D�8�_+7XUE;����zߋ� �Q��I��'נ�Bt-�F��0�����5s�i ��Ei^	�' #�u���?2!#N4B��� ����Rт���]�lԚ\7c�1�2ݝs����l�50u��������(�며*1
Ǥ��Ƕ����R�N� ]���ץ���3�=�;UͿ$��=UDH���{2�D�Y���@s�3cK�)�ޚU��q\l�U�L**�x�tɰPn�@*:�~g~���@ƍ9�]ߖ'�N�J���OR���m
�{�k�h�,1Fl��Ӫ�(^�@p$�[1a���O��꺋����8  ��3a�@�)`� �;�"š5���J{�YBy���.W���Q�� �� �7H�	����{��%Y�q>�ա�p-C���Vf��M372����c���$IQ�o�?-�N#��&?�*�U (�)�HU�!���Y��K�P�����+W�`�4�v��:)f���c���)f+��ų��[�����ֿ8������ GH��m�A�~�oh�J=��Tƺ�HQ9�qx��*0�=f�� �q����һE�K��Wݣ�3�;����A�g����N�ǛkGv��eڑ���.��>�Wv ��csU]Bm��66�X>d.��CI6_���ᤶ��E�P}�wW�˽k�³~���[���6t�1'�hdt3��2\�w:�=#�;�f!M����6ĴwHr��1QҤ���RN��^�s�4g 	���h�.�����Niaq%	���ΛCb����~�0�LBW�2ޖ�FG='Lt�(7~�YŦi�rY����H�03W�k�W�ȗ١�q���?΀�J�����BВ��$3�Wn����%�%��#}�7aɂ�

9ߩBdT���T�@��y�2��°�rC�ɓܫ�YwM��O���.�����>��;�uwl���c�m�@�~�C�6��O��e�T|��{zvO	"G�J�c�k��e��y���ʾ�z]���3b�X
6�y�d�U1}4��xA3�L��)��6�"��ӈV�u������'�[�vJL%���H/޽���~�	�����_���j���W�X����r�����I����R��)N�� ?�嗶�wE�Xijj&�8;~��츝�_��	�׌*�t5S��IAň�Y��%��g�灧�)6��6�����a-��Ihʰ{N*�P}�fé��S �$^�X*N�4Ͼ3+*&Qw�wH����9�]~m�UI���^�^��hs�x<�*��V����f��+X]�M��=ss���B���]tј�Qxߖ^�:��6��#׶+ۻ�t��"����
"}7��j,5�uj�)��4�IX�#(dJ�iHM����D("D���J�z�GCйӣ���`t<|
rm�fa�������e�Д~�>~���#�as����~�����J�5܏/����٩���\]�b���Y�VdLͪ�@��p21��Le����^.�w��kX&���]{N;�jO��2�~��uQ"�,d�̥]�Y�z!��s�+�k���Y0�>G��䇰Hg�
r�GO��	D�8�rӉ�>	��)%QGCs����L���OFƄ����쎎�F�r�ɠ��q4�[�*s�L=�1>�Td, �����c��{,8)�+�`���ˢ��B�4�&^��
����ER� �Bd �`lI&��}N�o5�`d�� )j�0�
}EiT3��TXb0�/�+h"���o���5���;膢��s�~�诖���y��]Ϸ���&F q���xJ��K�7I�[9V-*�kj4� ���XA���l?��6j��:5,QP��8�	�Rtz������?�����#ɑ�RVh��RF�:Y��U�L���ڮ�U�5�`M�b�G1��a���y<�};.�Uadd|�(�1�9��u���2���^|�\E�wIKsd��r.����c�f��^j^j^�Z��y&7�"���-���8w�k^�mnr�
>vw�^�A��z&	0Pl�����Ύd�
����΅7i�k���W��/����B�FX�%��8�	�r������ʾ��Q�97g!L�N���K��HCn���_���ԂS�g�����ժ��5҅oMw���q�IЅ�ݤ$�o�+�Y��G|���n~y���y�&=>l��u�a�qX�eS��[DF����� ��y՛Z�ń�݁ò�t�O錔2�����}T<�����}�-~�5?��J�����ۜ�{���]Zs�h��
�=�!�nC��b�Q��{��#Ǜ�q<���{��	��МcE��Mk|λ*�M�]��HL���+a�`|���Ց�oǟL~z^<��*���_��x�d������&B�5Y�,rΔ�aa(��`���@"�e�%��Zj9�/�0BTl�YH��Q|���Q�Dz�-�/H�H���2&Y���ޥʂm O��|�����%՗2���Q����e
J3U����$f�r��+�[��j�dZ�����±u!���K��ל��Kې��*v���ZMRϗB��d"�~�f��!�%�OL{���q���6�7���b�뫍*w-����6�{6ͬ�2�h�grE.�$NT�8z��*4�VؙHxՏ�^=3('���8�����|O@��P�Ii���Li���/6�����yX�5n��穭;;�ߙ�=nƤ�$��VC����
.Ha���}qm�>YY�B�ьa�*�c�*�l�~��+_m.� �F0e�QsQ�ܑ��9z6���6S[@��&�e�\�k	`t�?��8w��2"�/f���-�?���N�xqX9��eh��!���ú^�&���FQimy\R���ɳ݋�c2֯�_�N��캅qKl��¹��Ih��]5����#�<�x�{�����q�7.��ܙ�����+�#S�!�,��)13�,�D<ga�f$ ���'gV�7
,���}5 �7�7�O{{� ��6���+�Ev�}��� Zĝ������M���C ��n?+���Xk7C����}��K���v|�	�|���]X�������׊>�ٟ~���A����	��=���<A�(�U�p��=D��*��P(�� �5$�����? �����)���T�ze?��J�aJ�	�-h��ע㨹,G�-��i�M�ek��yѶ @�u�_��6icu�SS��Qgk˂\���^�JE�i�7�vX��B[��
P�+jҒ�VTĉ���ұ1���D���H4%��p,ޢp�x�fƮ?6��������&�����Z�6�>� ����u<V
�x	�p���D3��%�/'S^�u�םD]�4��'
�,5�[}]�ݓR�HΔB�O'�`L1|ڡ�6��A-(!�<`{x��x����9˩M�k%*�_�;X��i�hRB'��@d<�Bq��55������A3��d�)bv���iY��0�3p�&��x{�z�c
���/���!Y6������4Y��*��yL\\��ͯ`����rz�8��RNڬ��y}�d�\�	��A�Zu	'.ɯH�E�ڄ�] ��o��A�,!� ��|�d1o=������i0�ݦ��d��F�v��PF=ƻ���ơ	�	|/�ҏ�^�wGWRX4�I��;|n�z����H��o,�虙�3��sF'y2���'Ym Z}Ecܞ��5`AK/���3��/�C�6(�XS��hȔV"z�g(��I9_�,#͠���� 2P>�7f`�4���	�P2e�O !�y̖���tbcS��;������?�Mu����}���W7��T��e3'��fC�~��"c���<>=� �֡0��0���g�dp#�!��eG�F%'zڒG���#��C�$`b���P����~� R�k�������(����ռ��G�j�C��^����-v���zOSᝒ��
��3Ut27�q.��s�/�b�K��n,�o=�ъb�N�UC�77��wnH�l~2�\��P��A5OK���fp���`Z
@%,1"@r�0�����1ӏ^�;l0��!��{M|��B�X`{Q:��'e�aI���L�=K��ᾰL�T�ޥpXD}k�ZN��km��O��E�Q7�&H@'?L"�Z��{9�j`��"�0~Av��7^7��Yp��/� KjV8}�����J�<�5!���@L�6���$�\V�y&@�(�{���"E=Q�Tn���x{��*�~���]ޗ/�3�.m2�`,�֛��kM'cQ��a  ��)�	��>�2�����m��u�M�B�wg�<��Eͅ�'�� �7�B]&*Z853d1��a��zS�-ab��/�� �T?�1p�C( 4�\�B��
����.XHb�r�! ���x�W)���R�3nL��>���y�c*����cQ6w��x��7��V�T���Px��,��_���.�3o�� � ރ,R�`~�46��k��):� ����7�+� v���6�H���6|/`��X8w�( { �;B�p������Ml<-M��Ƶ-"z�O�S�K��|ARar6�9�[��+;��u���eu)����7z����I��ߚ���Z4�S*�=�a.Ҿ��á��w-5�(����P�5�܀X���Z��Anhb>4�qR$b�}�����њ ��h� `��A�����fkkkLu�B�N�F�p EX�1�R�߳�=2e�á�#��񼤭B@h� �� P��nR�TEក��]DFo��*x��%Ȥ�dd��������	��%%�j62K5���J.Q8�t�v��W�"�� ��)B�E���������hݨky��+�)2V���%|P�p��Gi#1�%�1N�E����u�_����M�zk׶d��
����ۊ{v��ȴ�ʦ�����~[�6%�'Q`SL/I?����u�h�������@J�Mw��֕�[JHL�o�	aڅ��L0͂�����6F(d���`��4qb!2�X��T{�d: ;�����.Rw�!r������rH�lC� �ٳ�(�:;r�L8\�U���ys�cw��=Uki���]�){M\c���PR�>�a���û�&e:�&��� ����W�p��rGMf*2�л��b�Z GQ?���|�S�)(��#K,����l&w�B��8J��c��s�������Ƃ�Y\�=�7�������4x[�28Tș�ၣ�)6`s	r����[�GPU5��<q�E���1�D�L-����4�h�w��?7]7�ܖ��UU0<@��dy�ٯ01H�$��Eh#�k0ICS�����.�ۜ?�ؕc�T��Ik�[�eՊp1	�o7�O��H�9 1Hd�6��w
$Hΐ&f���X*�%�����\jj���(�z&��Щ]�-�z֖/��[��}�)Jឡ&t�� $Nd۾����D��)>�~�iݏL�	#�n�*�H+�ī�#�hA2�0�sy�q�0���_����XʉC�f%�'�}���[�)�f�(OA�������_ݎw�����4@\?m���#&�̺|�+2t����K�k��
@���=^�MΟ��dUd���"}��z-�`ȓ�����#��.��;j��r1/s��/{涱������0t�"n�#y�K��1�?D`]���kW� �~]]���ԧJ:���0<ssF��+�m�K_�n!̖�����y�[��q3����'٥>%�$�R<I���@��6�r�L�"�T%إL`�%W-��FۦE����p��!���K�9���TVJ�+:�珙�'=r�=e�+�+���=�r���u���c')H?���V��P3�)�8|�MU�ϐ)�i�ه�T~���љ�>�����F� ���	L�����cVϊ�u�fo=T�����7 �}���yu'�:�&�
9�Ҷ�u!�v���2��!����v�)�ga�E��GJ)���c����W�m�GNs�Sg������" ��6�����l�[׬��O�q���{��9�
�0��-���2hZ��A@�Vc�眻ٺ�W���?${=��|~.�va�<�5L��M�X����o8�Qٰ��p^��y�R�����^�F��}h�CG���XCpS�bIk����A��[��N�7P����(�2�\^�+sF;�`��d*����>l�f��n�B9�\?�Bh#f�s���EO�ܙ\���Q?���A�����cG���p��'�����bG���uiY���t�\'�
�~����^���^�ļ�t���B�e�,>q��g��dnp^q��ږP���G���R��,D����B$�P�E2fM�H�Wz�ԝ�U�dq;������7��p�� �^C�t6l݁�֑bj3�i� ���?�v!���$�!����+\Ε��'q3q�nm-������ہ���T(�nl����D��3g����?"���e���d�E�F���~T���V�h�s�.�LkYǍq�P)*�� Xh���"0��)v%^�����.�_��K��I/��ޕ����L��h�KUs?�B�UHG�̩Ĕ�n�b��*�sw����&��9*k[α�
��M4k�c���?�B������r�-�:6|���
x�#W�b�M�+��?�|V~�%[3~60�:ǂf�BՙP2A�C9�ؿ�:ֶ�kJ��I�N
�3z1K�l�|�0@h=��7�*�?�M|`���dİ]':l9=:C�UB���^��Z�;�w��.8 &<�^8@�$��N���R���å?fh}a�ѫ�2�ޓ̠�O[�\ꆵ��sc��؉���L�Y�M
������6�#��l���1!�t�j�<��#��� a�ݐur#3=�
m� �~n�k%`���Ч�DO�;3]���h¨� �d��t��Ġ#Ŝ8���c����s��S��}����ySha|��_��-�A��SR'�cG�a���d���P�kLq���I�H���,:���Y�tyI�ї�cXl~ێ���$�(�Y���6}+�z�r��d�HF�{'z�1�}\���v���v��0��fU9g�D�JJ�G�u�ˀ�4,X���xn�q )�
h@4�� %@ڿ���?<�:�\QWל9Sux��Aɦ�R(lp�����Ξ�`%T��Q(���rAA:so�`�ȉP�PGUU�A�B�"Y%�7sv�2��O����Ŭ��LѭF�RE����gϱ��Q$@�&�낝61�������4,3��z�r�-��t��2OS��k-چ��'0�����`XS�O)�"��Bfߤ�a�[���#���o7 j-X\�
N7��3P{_}}���퍍�cm>_�* LLQ@TRDK��/i@��".ʐ2D @�X����������f��~<����n"����h�W悇�d��pz�h�����,Yj�KG�����p���� ��t�0�a"{��R��c�=HBcR
g���2s�ݡ��*?״��
��3���	R�B��hYP���,n��Z���Vs�e3_�����sr
�d&V@��~���w̌Ү��[�`�_�M��״i������0G�h�(n��jG#����D0�2�n�l�����;e�w�M ����s�ΡP��Y�2(v��7�k�u�7&珷�:�:!�0���B�X�    IDAT�(sg� �a�+��0�v� �p�TD�=�����`�Tڰ\L�������X϶�a:��J��3@�r%��@i(��9�T�d�\���U��8� I�X�52XS}���l �q��Lٙ�;�7��;.,?_���7��ܳ_E����ݝ�$��F݋A��3b�PG������B��ʧR�&���]�03�<�����~z]�F!���9��
`�s;��`x�03�̡ ��3�	�{���2�ך�q.����o+�+���m��wo]�L�#2���p�
��&�o�G�Q��d�aբ}E뫝��Q@h��m�|��o>_��3�t�YXV�CE�'˪�s�6�Ɵ\Q��ެ�W����_�r����I 1��bE�v�ߴ�L��ǛuR�LƐ����xUp�*Ċ�j0F�f��Dڈ�D�Ґh��im���Rs�6�t���ֻ��:��]�w�]:�쒦K�G�?z��<_���u������%"/?��y����� ��0���&'��T��L2�:�A�W�4�O`�������'�> �B\�
s�A8kU��`K��qeEd>��/V������55nC�\{{��f�͵�3a��h�C 
Y/����Ӄ=�?)��:���KQgXvƄ�GK'::.\�p��^k��Z)x\,���k�r�%�|�x1�.Hē�� �wu �����"j9�Mj����|'L�U� �� [��������9r���0i^p�S�ƚ����PX�3�Ժ��~�TzRj�f�}5�+3����n�L������hC5�� >G������^`��	� ���@׽������
y$�Z>�W:Ҳ�"��O���]y�ղ �� a��ϣW��R���G����_ ����Uv�P���	�}+�
=��{��s e��n����D�5as��.k� ����B����K(�̊%�p�= �_(�95�0����/矷��k�͇7Í����|�5w^���p�����H��e���7��s˩�{X��f���@{����� ,�|� �*;a��\�N�@@LM�ck@Z��½i���?��`$ .���&,���ĝ?�d�����W�ò�vI�˯1O9��8R���# $ZU�"��f&X�����{x9w}��Zp��f�g�?2A0窫K �ٮ>(�ܾ�@� |��Z.M?Ć ��
"X ˧�R��C��Q R`�T���:��GN>P��c�mGp' �-)�?����Y��Y�G'6����C�p5��-o���#v:?1.+�D�'p<)1V��@��wg���F���O/ݽ����K_�	�����u"�DFϕ3=��i,��������Oe��R���*�g䢧S��.�X�g�y�`
�8���ج����c$8�h�D(�f��9�U! a 7N?����8"#!1`��@���2*R�2�?Щ<a�h��nA������1gʂ^����h����Ǵl�8�_�U��{4v�kx�(�`�� �Y_Z�?:�Zݜ� ���5;��@hb�oF�]��I^)���/MOo� "�RS��Zr�^ GǦ�j�p:3�G�>��)���y[�I�!D���8�9t(=��L���ax�F��Dy�����.g���iP'���r��E��<�OP�D�8�����1�#��/(���rX�дh#�� %fe{�t���+�-�uD����E.�R���2 F���یD<��B�:�� 
�NL
�U�����z�ܔ<�>P	�ᕯ�N{9��:bH�ׄ&]�cq9
��s��Ŝdڭ���%���!�m�s�H��F��~Z:q�@}>�P�
�"ǣ���}���������{zj���/k7hdT8g�S�ӷN�Q &�A�A���-��"�=�A��'�mC�e����k7 �o����@>m�`PX�
��*[z�+�	���C"�bb���DT�lT���0�1�S�,�W�Ϩ�u9����9��]"����NyG��duW**��.���H��|� $F��z�� \�M���ʌ��Ah,(<��bܤ�c�*UQ��'��aj�l�4��>.G����w##"@ˏx ����{�c#�[�4�r��\.,���n=_Li�f�����KH�����b*�lR+��}��@2�ӆ��<�T����g�v�a�.��u����B��� �c@� ���S��/?���_<�ga��|����Ȑ�R�
��8��S_��僃%��i�钕�J���I��V �G$2aɶp��94�~�Xy60��ܓR�w�<��x����Eu2gNB�)�����A�6�?g��\�����o �j��^]��D�6$\���S�A����]n�_A������,�ĵ2>�
��Z���"D�����D9 r�I�< 1����/���߁�����^��D3�3���]Zz�7D#i�����7�-nep�{�i���Z�TX�m���d������uu=Nx���t�s #sF�v �D�H��H�9L"� &�S���PTǃ\�q=�V�]�󩫳�`�YR���(̱�O`���4�ϱ�s��p_o�{�2���#���5�ML�r���Fq�غ���~��o��v�d���|�������|;����; H!ө�n��
��a �����'k�� x�/@�=��~��D�w��L�L��N!���}<�������,9�@�A ���A�,$��ˬWS�e!�kU����찪��jh�_�?�6.��>����x8�´,��&�7^6Z��м�f���u��3C��۰x�v�̙�))�춥я��������������)�A#�H�B��D�ӑ�ޒ;�kp��]<`$�Ց���kcA�Rwcؗ$�#����F�gU��+�~�O���=��<��D�V�Ѐ�@1m*U0<J���XR�yX�PHi�[�Th)"iR��P��I��ca�Utd�A���J�(wv'���l���wo��Lf&�M8)��M�(��{�9����#\������t��P4�tI�T3���:����@�P��$� ���d����R�8&�w���͌�� ̠!����D2Ύ�������w��<�>�������1�bn/ �_���~����D<tδX�	h�����G�,S��dB�F����W��nT�{�n I�Q 7m�R1xg�36�u*�xn�ÎfK�&Aiiu���ʛ ��	%�XLǋ5�~�Q� �0��zMq��娺���  ^�M ���>�0���nbM���c�,Z.�RH�2��jMqmm�`����w�����|�O'��^8��-���Qw��mMJ�� ��� 2R��$6͍�H�~� ��_	Vn]�6���ӆ����~�qr���0��tsU��D6	�@4	F �~�б֊_.��c��b��.��D"*]Ks��y;=9a,�ș^��ښ̮>���KߪP�������r���mȣ����U<O�]f�M�&�N(�}���CeQ�CQ��G�-�um��xI����*�q
r�x�,O v���Ή3?H��i�^�0�K��r��\�]���k�SUs�t��> �u�8�}c\y>��[U�}��@��^f���+K"��!�!�˲퇀�_Y��� �8Ta� T�O�"B�,w��]Q ��16�o�3�����3�/�����>6?]f ڶ'  Y�	
B���s�U3[ O�V���|
/���@��iy�c��%u%�L��M���#{F��i$G��'�H3�ݏ`W�d f�]*�,��s�̹�,�3q�i\9����ȧ2�ʤit�����IT��)�KѨ_���6������
����Δ[�.j> �ѵ����ܨ�Y/3C�;��VKA����W>�_��Y]�����)^ �c�_4KCd�rd�
m`�slkJ� ���	�`0"��@�~�r$�\PR��(��Q�Sܑ�*��$!���nHj�M�����������:@�:�P:t�%-((ȡ /2�����
�����Y�EwSO�(8Q��StE?O+���g䬈���cxxa��䚀�L�]\[\[�Jr������:r86����o�I@5�-TD{�<��\�o�9�Ս�K��"'��7���}�L`��E_�l�XXB�&�mqej�bQN=7�h�\`����h�e�SՓkK��9���{�UM% ��D<�� ���+x]}�!���cqd2��X�����R�Db�H$Pj��f��k%ny�Od_�<��ۅ����m �s���;��HȜ;��Hs�1�	��=X%�_b@`3�U�/���K��q�,�����@??�s�g`QD0=�\ZZ��O��W �����0����F�����i<�'��/=l�ȟ0�J�6����:V��HBZ,i��C�߭�m�5�0�y0�c�2R�1�.݆|鞀0X��St������p�ᣳ���h{��K�����fy�������A��C��ζ%ѦB&dޕ��#�CW����䩙��+OG%��;�e��t.�d��y`uu�;(H=i�L!�p0����+�)
@�o�jfͶ��0*d�9Ǻ��� B�m h}��ܰ4�C�z��C�re���\}'__V�]�|��9���������%-88�ˍK��Zzh.��q�,�"�+�
�����t�s�����0�qJ��p�tC���f�is
bJ�����ti���b562��`��G2����6���|R�<����L�3ǰv��o��27�(icj-���:ٟ���Ď��Ύp��������*�Emh����X[4-��31�H��x��'��c�!�y��%��CU/�������?���H{��\�`�ټ  �'_$#�ȩW��$��lY�E!� I	��ImT��Ѷ B?� �"��[ ¦3�{bp���2�yk%��v4r�(���͹z �=�����o�DF֣ K�H����*5�Zxl�e�
C�������)��O�����n��@X.�0�@L~ݳ�+��,�Hkx �;\��c�T�@�����
k5��;��K�7�(����̪�4�_H�Z��?S��U�Uk1  ��O;���ixx�%]����s��lXF��sTG��ǏGGÞ.&�{Ӌ+����	�mw�|*�Z�[�
�'%�O�)����ox�&��ϭ V^��
0$��d�<��Evp:(4�^dg���3'e���D�Wίh�
Q���c��G�v�܀tܚËքRY�R�ᔦ��Gpr�e�Tb�!=��P{��� 2��\Ehz�sᯣ��n	�K�+�K����
 i+z��0�����_~hZ7��Lt�,�n�����I��K�/���F�۳�+Z#�°���H� 3���`
��O�����i6�	�xw�<V����s�i:��8��Rт5�bҩ�ڴ"�CZ�J
�Z��Z�D]�@[���Gk&ٲK�i��t������c^"@�dyH�HP�.Y��1���=��Z
��lL�٣�������s���s�g���[wl�:��������=���Mϗ�\�nąe>E]s~�oΧ�[Z¿YL��F�(@�#�|V���;xzT�(B���ZW�S���Ȳ<���z�R#¸ȇ]9���͙��������C0x��>
�������v~a��q9��'aˎ�!�o�>�&�EU��b���!�D�f��H����|��C�.R��Ij�oU ~�&׺���:�Dn��\�! n�D .��ܼ9u����G-r>O'~̂�r�Y�JK���I��Y��u0�r��p!�M%9��P���a���$��=�_���b��3ʻ����7����ʒ"Y�k�q��(>?#E��Y�m�u���}������~6�2J�8���%��XeLq��"�꾵p���[��,>km��T�3#��` c�2Z�	#�bc���K�}y��Wn"'�>膳���z��> �/�oj��?�B��6�5` ���$FE9�I(�����s��I !��.��P����dŠ��:�`Z�5t�ZT��1A ��S޾��ꙝp�OuM��݃�w{��3`������L���(��e�8'K����:z+�~�1q[{�uo/���/
ks�:Gu���p蜐`X�2��b�8������2��b' .ݶ���l��K6� �M�HZ���. ��xX�����_>m �Y�X���lZ������,D �2��Eܼ���4hX� w�}]^n�M#91=<��(�\�@L�o~������Ąm����v��6�I<U�X��ɔ��_;OP_��e�gl���((��}Y11��ܘ߅�����T6[DV>;@ �2�|����On7ߙ�����~r�
��|��v%h���½��JiP����ȧm.1g��[�uT뽣M(�j0��N�SA���t���By�a�` ,)%���X�]@Qj
� ��� ���y�F��D��Z-�3~@������ݏ.o޼雙�����#��ف���'+(-8 ��y/�)�"��w!����Xh����O�~����X,����������6}���	�R��?I�+:���-5�ٻ�'0Ժ����e�X��],�2�*C�,oƀ�1zKI^��'Baz�b�E%2�qi �A$�g0@g�`��(��#��e2%(1�AI)���dr��*�J����jm&KM����QS]�Y�<:Z_W�px��`��֡3$^���`P)F�� Ah�
K<��Ѱ"�Koff����F��u���������G?�= ���]�b��%�1�.���z��
�FY�ڬ�w��]�rgE���ᅋg�.��+�k�θX.�>���v�j�]{״�}W�Qh�Wq�����C �t�(�Q�@R�����D2; ��3�oj��2��o3H	�R)%����~�~?���/�*�q��>�����#�yf3������*3g�2l���H�*ZY&��19qF�H!�� ��
Q��יt&S�I�k�Y`\���(SK��*�(Ѵ�c4�/��l5A]2�%p�#I��U賑����Iaz���:��ТE�vt�h���)Il��H�pR�c�}ʚ��F |]�y%'��?���8 ���"�L%B�

��u���̹ܠtz��K}?��T�����A���ש_��s��������Z�/?�}M}6@ ������� ��� �ǧ�_Y�0*W�8<\�@ 0Yc��5f�?9�,�	�x�;?v� `��x<�Nz���T���Xrr�2Ԅ��2���glf���#���� +��B�l��%��J(Unm�|��7g����%[ƿz�1����S�O�#S�~��AT����_	����S�-�%_U���r����
�^(���"n,0rCcW�vAlƋ�`�~��x>P�
?�H�0}��[� 8��Uo�N��_�5V7�+��K��=��4��aJU����԰��+����[5�s`�Q�� wqp3z���t��L�� H�U�p�hDJ[�@�H,��E�"�[�z:���Hv��{x�LNtd�5;)2<<2��m8�>y=�g}<ts�š#�`�L�\n���"��w�~���'O;�:��*@@nՙAl!'l��V �޳8��~��ǹi�!�)x���Ν��Z�[+$~3b�N��� `m�VK �+���bmAٶPh�]G�o'M>��;����LvW����ɓ��B�@�z��p��<�W7��'q��Տ��1��
x�����>�� ݸ���+���7k4|�_�7�����`�X�2�C��bj��sp���i4�����K:緢;���G�{��\�˷oy����/���gx������?�j-T�k&�BQ��X�k�>�Db��۫�ȽJ<�?44��� ����a�22��G#����[<�swC����M���|� ��u-<��BЭ����Qt�.vܼ��������m��=�y��w��VP *)ϵΉ�SC-9vE�]��#�\l��|����'    IDAT�ԝPSW�u����2$	i	""�P��h"D����Y�!����Ba"�C�.�<L�A�H}����[�Qcw4+�R�ngϹ77�Aе����\����|�����w@�Kz����P�x�������
�x_
e,�%3a�����k/FF�M�1���#�3v;�z��GG���G_<���h`
?b�8�e��J��VY�*�2A�ө+aM	4��E�>�vUJ `ϫ���b��!�Z�b��� �]1uT�����\~3��D/	/D��2����9�K�����X��L�0k�S�a߻f_}ssscnA�|sЊ�f K��� �V�("����m�,������в, }p�+T�'�X �)�3i �x�A� �y�ƃc;���1h�t���|�t6�mx�`�g��A"1�>6�z	�/��Q�q��@�y϶��׫�Uق�A��u@�۴�J�fzWu��8�[�t�sce����v�d�ƹ�ۿ���ڎ��!��68�KI��# � �W@��BrA5��.��
{�MWh����8�&8�|�3�!�D,�+�p7�hdёڎ�P4�,V̹�pt�� ��<^=t�֒�X�>@_�o���Y�m� @�n�Ϯ�\��ɳǏ���a��0H�ҳz���f��|6���(el�D�w�7����K����J .[BWJJè�ٯ�B?�\��)�rs�sT�����b�bowWW���:�J}�bAHV[��q N p�6�����`40�DhG�����`8��	��!3mV��فf}'bC6��#Tr��2�`݄���9/����T�!�= \�'�Y��jҩ7&4mQ��A 9)�0�s�/���{K�}�#|�����'S|��x�s�@�Q(~�{���/�<�Ӡd�T�G.����"6WI��\)�J�E������|:� Ą���L�Qb6���Iϙ/BERҍ;��ٮ�m��.����q_�s�r�r��3��ն�&5�X�ٷ� X�S�2�~���rf4K��xQ��a��(k��χ,�焅��Tn���>*��R�\�m�V�F��&/@��^���L3��� ��>xx����WeeeYY�C3!���Z*
�i�H"/����,!)$ph��r|9��a��p� O��;�l��/F�%"�H�B�E":]������}A��GG����rwQ �?}U}9"�"l{e߽z7�����&��0q��hx��Rs��3d��-%W�� ��
_ ��,�G�h��)�Z�Sg�E�k����>`���̈��]�,Q��6�_�p�<''Y�|��5�<��	�u���u�]�w���DHY,�.%��, �5�L�pѴ���.��,sO-8�;�&�$��,�A�	��ّ�?� �"R�ǅ�B.�n'���K��~ͺ3)S�vHw��C���e@P��,�[_l�/�ơ �b��Ō�u����JੈD
���<A�;���F��o���+f�˲���܄��î7��'�lZ/�@- :j��y�7���8[5[�� � ��ФV麢.����Xvv�~CQ ��H=}ķv4+ )�O��(�B��+%��K���9?<-@h�,���������z� h���S}"�T��v��~WIooUUgKb^aH@�ֶ���'s�{k���m,hQ�!�e�w���o��ۢ���h�*��q9��9�^`����1��%B̀�T7�MA46�S��P�I�[|V�'����M �|cwU��W��zwZ�:����_�Z��QC�N�� �� ���C g�{j���@@&XT"����$�aX@&t�f���>� ~���z@�D� dC8VW�Mʔ��t�fB�Z�٪;/K.��u����u�O���<O&K��6oZguO��]�8Q�ӑ���7���ӞMa Iq9N960���V iP�K��O� �o���Ҙ���W�(�m^�3��f�D�����&����5�a���[:K�\Pe��L��(V�����2��E$j�pB i�_&J >l�������@�������w�s?��ӧ�z>�@�xk	�"��x��j��XNff��C �Ѣ��M%�Wd�<��k�F���V�j�ݼr�Vq�yA�.����l��<�� Ȁ ��*�6���� &�D�~��0�?��4����������sL%o���T{���U�!�����ߜ� �Y����NW�*�d ���O����m�e��r2�0Zo��ဆ��`�Y(���@�2'��e��d�@�	@aX��~)���}s����:��ê~�,����u�k;8��nN� �� ���Na�- � �2�$A#CD��Ǎ/��|��`�k��s�eT.�0�� �cz� w3щ= A{���& Qx5�LW���l��ז� @�Q���X@��� ����
��?�� �������1� ]p ���n��:uGBB�Ѫ�h��������5����w	t�/:���ځPo�L  i����-23�?�4_[�� d�����<��::�r�m@ �����ش7���w�7$���~"�����kLSi�d+Z�n�4Ж4d)
�PZ6��nK/Ci�`ai���HgR�@��� #-BYd�_*�Tu��D��:��8��wgYg3��=純K����8<��������������e�S@x��P�`;:��^� (@��
`OgN��Yp�*�
�X�CY���JX���ڢJE ���x��2Ce]������f�����G����Ɓ�J���R)-�J;|d��5����A��m����&`;��|����?���e�����8Od��3��)E(�.���}�����~IJ�}�B �'����f�`c �k $�(��Q ��j���n�iD����0��0��E���Z�]T�x���T<����ϊ��<�����vٓ�5�
!7� ����c�w�5�zf� =`�6�B s{o�*dErEM��T)�����b�ړ/�}tE$��0..n��U
h�9�~[�2U)*@�Ϧ�z�F�?��dVp�yԱ��Nuiuk3�9ޓv�?Ι�煌8�(>�󕇮RG�kF LJ�~[ ~��� ��������!O�B�1 M��I��b�yb�b��K��ۊء�����~�B�F
踕L���D���0�`h�ܰ48��@�? �|%����A����JG |����\��k�4>uJ��ڪ�?r�$����x�xg_� w�x�����s� �PqB����#�����: Wރ�_3}��T�/�̡�F��|}���9����32N���XY��s�ñ�]�q>n~1QCd�L@����Ə�$JL�,ۦuK��: C�o�D���v�?k�ź��
Jt:��B����!��a6�\���<&1Q���Oǌg�1���+cu��xVƥ����8/<H�P�:B�u��z*w��T����C}	�v��� z�w�t�&��ݯ�CxЙ���[��	<x����	 4��P΄sF���	�����d �=����a���>�d�ġ!)&��M�@A]!�.j/ѕ����G��i �HF�:A l�����WGc��|���P��ڥkL5�v��y]z�ӒiLfr�hV��g'OMyT10�� <�������5��۱��'8;�Jl�"y A-��mj2 e*�p��<�+J=�= c�����J�~�f@��#K��;��뷷�F T� v�W�!H,��[��E|iA�� ,��#�[^^&Z��2 ��@�P�E�9�fuj��?;�OCO���3ɩ�L&ϋ@;|�v�:c��\Qܕ�� ��p@��[<	��>�ǆ�)��4���4�C��
�5�:��I*:+l�~����������q۶� ��(!Kzb��ޖ�E7��nd�9_/ݴ(��V-�  �)L�S�J�^�P��?��:�u	^|1�� ���j5EM���<q����D%d��=>F�����2R:�Zv��.�o�'*j=gk�j@��� ��p���'>��@�M�;ޓ������zC�%uRl��`l���bH�$�{��tF��{��� �kFe`����;?������x��a�$>+w�"�2�$@ �ؓ��dE� �@�.���o��� ����v��^�Sb}D:ѶsU����	���P��`O��Wŕ��aFS\K���Q*�T)��#�������^����=������y�iDp��r���W6��qO �s��b�����/���z����$�TgE�J��R��\6�:�#��"���ډ�G5l��ߐ�Ƥ{o�n)���Y������50����5�De;Ȃ5 u��R�k�$h��z ��yA������������U�����6?^]++/䈓:{{n?�}���������eO�	o ���Eg��p�`���0}@k*�����Ǌ+��������Ɋ�R��~������>��W��*JG ��&	8��������t�tܻ��o*O�v�(�Av6�*���HIɆ7%�� D �`���`�H�~YGm��u@u��B"�[ִ+ET������偁���r���p�L��4];]��Lr�8��
�"��^�]�-���3�v��ߒ3�Vz���U�}�&��Oã�� �6��/���X��Bmn�L@�` ��;�
���T�������Ĳ�*6� ��/�}wLҟ���*L@$�2#G���q{��>�j�6�'\ܳ�U Z�Z��7����@��t%z|i��^�\�T���U
xKX� ]5N��t�ܤ|!�*~����o�ɾξ6����m��l�e��
�jV�80��ڂ ��m����3�ޭ�z�ab�%B�o���)� 88Q�R�c�ry���]q��Q�`!u#�G~3,ٻ�v,�S:����ؔ��N�#Y�l��c&���F��+�&s�} D�M7��ܠ~���J�H k/v\�۩D�H4�^R3 ��N��\z}�F/��X �%��|�M�=Q���n	Ł���`��R5q�rn�j���"��\;��#�ɏ�9�*y�"*�^�B�6�nY��'��A��ѿ��sF���r�FG�]�E�:̘'����%������8Ρe�t����2�ǊnbR~$�K 1$ĮI���+x�J0ޖt4��4�$�3�g�WA��8A�pEXT�s��s��n����<OB�n���m�!yx��{�����~�J��_��g�0%iYA��*� ���>7�2����"LPP�ڐ�8V�:T" @�0��Cc!�!�Q(�jZ�ʑb#��E�4i�01pkf�K-L�������N_̜�5�tv;�C���C��2����K�7�0:�]��,:�ݎ�����$��<���8�����^�ތ�q��[s�~ "߄�tI��f��̔J�Z�$!�Z%�TU��*���4��L�I���ˊg��կ��t��$WW��uF(�6f�͙��ޢH8C ��X h�-`}�I�7�?��r (<��7����A ���m�P�2�$ ��C�##�B��̔�N@l�r��M���I~Eo	������顡��!D ��;����n���;q����ͮX\\<Z�dw�\ބ�����8п}�# �)���t6;BwtqQ��� ���o�'�*�vs�U��ۓc�rE�f�@J�	����Vk�h0�K�T����� P=�BIJ��I�X�I��څ�����`��'O�,<� �U2)(#�J�����(-r !��_�����I P��"�7	ćԼ��(��ԉp s*�b1
��^��@DَW������X9S�Yy�oWy���$Gm�i��C���ZI����wk�/�+����/�uf��0D)[�y�i|��%X�с�|��&�''���n�ۊ��#�9������P�,���Cp4�� J��(��s�//N��M������,�=ss&�H�>���!�Ǯ�6 _Z�pa�W=�9�u��33(������l}��>�ih��W�� ���{䏘����G���@ ����ݰ�XY!1��^�rq"� �XP��?�;#HM���
��M%�>� R�����վ��(24�DE��67���*�L"!Q�?|��]ɘvu���B���4sLd�+R����S����w�cI�N�[<����t~�ُ�J�0��O&�.£�rX�NO���9�͍\a�P�dL5g��mna��ݽ0w���_k�N��;t]Q@m�^S�e�����x�V�@ vw��F
��Q(�����G	&&�kwN�����ǎIh�$�qF��c���L���'�w�酞n|z�{�}B���7)�{R �6r���F_0 C �? r��111��� ���PK�����Y���J](�X|u�T�g��ݚ���ְ�Ɣ�QĖP1�G�@`s�� �pUm��L�nzgm?�;~~	�O˖�u�#X��+G����b�����,PV
c�~T0̴?�,/�!N���g ��y@1��cuOg��s���{�����nN�l�c�0(��?�Ԗ>�@�T5��g�J����1ه���??�$�K?��
m�tX�
��Z"�-�[nO���z���53��|�I�7��h"����B�,%/��i��m��R6�P�a�M�t?
��i���K�P�����b?{���\�53K�UU����/$�z�`��,ZH����c�xP` y� �"�,:V�u}0�������^�ډ}��t���'Qm�#p���(��t˭f��(0s�n��*�r(��p�<A���`��3m�V|+��	 a$�R�g2��?3hf��gY)�T��}�@�$E���6h�
�O��y��A���rqKF�}���w1�����������Ƿ���_x _�Bi�Z��_
�8���z���T����4u�b)����+W�����!#^I�!5���RZ���c �:;��-�Q8aSwV��PX�����7�"��o;RZֱcG�5���}������>�����;k�챋''� ӈ͸|6���B�b�U���*�,Ҋ������׉D�	�H���i }@����{���@�;8� �k�f��m�ם�3�$#�ǗH$��D.P/��c��٭�@X�_��������X,�_,�{�����{�N"�Q�u��� ��g]��z�$ڒ���9SrI<���l[
fБ��ս�i�Q�Sׄ����4�V 1�*< G1� �)Ԯ�\�3�B��Nߴ�����Qo4�.Ghd &@ٿ0(7.m�O# m�Y�'���2���s��h�h�hK����}&��
 }����;�]�5�5/�k[�sO��g���!r���]F᰽��|Sy�͎2�z[���O��8-�۠�����Z����#
�*�~t�1��p��U��u���]�2L�3�Y�'�x �#��sD*Ua���x��?e�89ER)]R*P߾S`��$�@t>
�8r 1�7nqir��-����7�j��ƀ�2�dܗwn�:�{�i���4��s����moC�(l!��q=��;w�Y�.��ƚ��#��ȍ�gg����89�� ��/\���g�����~D!�����P�s��K�o�s޲���İM��|�����=�Y���{z��v��3�M�S� ���2v��kы�O�BKKnn������Aa�q `�i;��&�4�7!��q%����p@NP,q� ?�R)�W��WZ�u{�B��P3@�̕��C�����h]VW\T*p�a����xQ��~������{ߙ�P#��RB3!i���>���>*.J��?bzcտ�\*���횹�kז����;��o�DH/^�-    IDAT�i�Z��>;9�=p��\^:;�_��������?/�̱��d�	UU�o����R N�q�9�� ?F���E�wj�Í`(M ��;�XB�B�Ə��p�ޥ� �N��6�p; Hi��
�jb��(+6#�hI��T&1a"0\�"J
����hH ` �
 ���uE�����n���幙4Oa���f=�E� ��S�)S��	���Ԡb�(D\��U���v���m`س��/.�x'Hk�uu��g2c(y� ,\� ��6�^.�
ɐ��~K\F���t+���\��[���랚w�C��f���Hr(�ZDԧP#v�L��O<x��z<Q��}]��j�P�Z�{�w�S�N@ Gƒ< ��,A�r�滵���g���fD�@��J�$W�(-� ���������uya���=n�v�ff�0�G+��B h&��oR*X��*f��V��|^{^{�偳ݓ����=����r	��z{al�A��2���������8mf��eC��:�jFG!�ik ��Q�_�p��O�b����a%J*�@1�!��3G�7t�V�s�&\�3.R �P ��M���.���p���b�P�$n�HB�b*�	��`n�}���ӧ�~�N �s�NNn߇s�d��IjQ˥����sۏ��}u ��n��i S��� &�Q@�S���	������]ǃ��!���E�ؾw��}�G�A���0���vRw�ض����O(��£%%M*R��l����+8A�W��i �{;��buEEIv�_=����N�G����S��R���~�% ����N�%p=(0�DF>?�����W �ᅸs���ᅃ]�
����*�w<bkP�̈́�QE�H(���C�]p����X����ɀ#� @]iޓ����1J�X*\8���'IR.����pmd2��?��͛C'���̾}����QB����䎤��Y0;qs�#'7'�����x[���J0pMB�	�J_���ꑒ[#�`)/,P�@!��L�ImAH��2���i���ęw8j���������/�:��J�����@�r\#��.�����Ĝ���5�N�r����0l�����#�Y n�5�dP�Rv6f�����7��  ���\�:���Ԡ��E�r �GA��
1�8&ǹ�D��??���� �8�� ���J�m��n5v����Gr����0��mbRbS��.yމ'&���_�UsW���(:hӦ�M�b��;�i8�<2=*H*o�g$U��L�BWI@�q�ԅ*to��{�@!� ς�tt�2̉"",8�]����>�p4�_�Ȉ��Q R���a�?.+8p�Ieѣ�2�õ~~�NQtuQf(uײ"m5� ��=Ey��7��e��q)�z�n�+=��Y��e�ڀ �VG�(a6��f�Ӫ4+�A�G`�@� @��-���W��f�
����[��z.G�Vb��{��W7�k��)..>x�`O�N��{��֟�?#9c��j�f�c�M��1�+���%N��3Q%�N�IJ��f�N �;d�G�ͦPG':�j�M�B��JV@g��Qu�7_w��6�a��RE�@��x�
^��_:ȟ>���Y�,�� woqO���Ȃ�Y�w�̌�I��c�DAZH�Aj�N���.+��k��`l���﾿��W�Lie��v�����'ؾ��iڂ#,�M(U^�q}���H���ⵆ3Y����78Z��?_�:�a8 � �{��p���b�N=� ���Е�2�i�R�nqll�'K+�����a5Z�rj�8��h\�Ke)I�X6�|�*����7��/~G8�cx�V��N�2�%-��q�}�V��������C_=�(��
��7B||%�W����WG£���D�B���}에�-����Ԇ1�e��ۘ��CKJ�\�C�����(PH�z�r��
� �e���E��q������!A��y]��������K���xJ���cy<߳M��tJQJ,{/;����l�������?4�Ө͖-�,����/2 ���]8�]����$�$+�0uM`:�:����z��<=���q�AH�����?#OA5q�׾06i���VC ��Hl�B���҅9���'ԓc��.]�L����鎹᳕�������(KUH%�[��}�XL�ɋq%���75b^-F^q�?$haՆ�ԷېNH-T������4Y(�r���F�T��m��s�V��z���࿺0�C�rjy�(��RdK_��Ώ�y� GB���������+�`R�;v��e:f�����1^ן���'v	boǪT&lV�Gn��e	k� f�d��8�������i�N�8�KjwD�rW�.Hv�Z�C�Z�	�V݋-!�*�%��Py_x���b�}�v5P(m��o���Q�):�p!�1����=�H����޶Z��q;w�=$�MI�P>|����}��G�;���a jO��'RR
L�â���z��!˳W'���� oL5��Gz��� �N�U��86R8��&0���	Z�}l�������׋'n�~ ߠ�5Em��R�0�,έس�����]F?����� ��x��岢��
wG���N�u�������+�/`4]�z�p�cV��^�հn�5�ຖd�+���.�H���c� 8u֔��v�onu�ј�G���K'�|�9�cǥ`��m����k���}��cx���W�k�Ju$n���RL�4�s�x�D-n�=��0�p��1`�vU٦�T@�p��e�b���/�����#l�������N��-+��Z��۞o�:`Wo�~_�&(�@@cЪ��Z��d�;�¹G��\6��|�/h O�w�|��"@i-�%�+~�aϞ�qLC�B� �゘y\���o�	T"
,�⥷��qK��
p�7am������5��ܒ��c8%kI���{#�1��3 ���c�\Zk�hS�x� ��Թ�.�N����uA;}�]�����4؜@_�:yv➧ h,G[p�͎�*5�d^��!dE��M>��]q	p�׷�dO�x<�ya�I@�煢L,��,��Z3�T-��mْpp �'{z��EI������@ep�>A}���U�>6��*��~O�b��]���C 3����^J���^s>�V���Q��0Q�	 $P�T*��&<{��y��QZ;&nN���k� �� ������4��n<�!Q�����hRmr���xsĨ����p�y���qy��k������j��B��O�&��-�|�:�������Al%��A wٲ��	`>����o�p�^ �ޜ�J�P���3`��Vcڍ�=eCva�XI�_�r�؅L��*j*�
D��H��_HZ����
X�v�J|D�E�J�p��K8�o27֕�6655�mj�4� ���0Ώa,`D!%�g�C��
.��J�d
U�J�O���/�= ˉ��" LZ����X��eW;Gړ&/ �)�H$rT�#!I�4��UDD��0�d���TF�I�\.���x"�1,&#Y�(c� ���:��we� mQ�N��tU6\�D
B��� и5M7��{���	�0�55����
h�:�Q���ח���sc�b�����k�BUxp�>%�C�N���0W���B������f�C�2 ���! ��X#����|� ��U�H w�M����צ�:��v ��(A� �g��H�@].���jBQ��dƓ���CvuÅ� ��lN4W�J��� �h��	���`���wh E�
/� ��"!♜�e�����2�D���Q��C��2&���=�|z� ���0"p8���3O�������~�B
t��ޗ�W�1|,�� ���"T=T�-��Q�D��̻ �\�I�"fV����m�p����`��U��� ��c�Z# LIɸ9�}�������U�y/ó��6 �'H�Ih-�:/�D?�T�A;�A�ϻ�~���M[���f%�T�ܘd��ϙ��N�K��:r�'�B�(wD(��
U�Ӷ���s�-KM�I�9�L=K�����Y����5n孴Z
7��4*3�J�Y���3��w��Εqw�ݩ7|R�����;^�+����Ւ2�%@�H䔗��Ɵ��+�:"d��6@Vtlr�~#�@p
����9�?�'��q]~������� 	 <�K�X�d���2{�D,�}������mK�6�T���ۼrP�d���ϙh]���+���Nܻ6�m ������Oxd)))���D�cr�),��H�o�3�!�;���0�_�ڕZ����c�V�>��v�V��ȓ����DA��B��)��ql���S[Ց�=Ð�-a��>��
�LS�����vߞ���-V��A0NA7��3P*�T��'�0��t���s4�4�낯���Pow�Ⅿ���se�O��ryAN���;p���4�4�y�a2*|��*�l���Y�\N����An�Z�&��ws\n��͎�卛qdpb�b%�=�&�l��$�����~�$GZ�*����X�������}�K��%��� @��r������%���� �zou� �ҵ))�s�|����*�R�k���E�pl6�	���`3��/��q��RO�O <0��1c�p8��6��H�B� <����i��)�􃾁6'A�Va,S(Z
���q2c��nt�^��3��A���B .� v<�xʽ{wÿ�;��4�;�w]�u%Z�fKV��.G��y�"�6�=((\S����c,��[u��hk,������N�(uZ���V<����.5m\���\���-޵��v�6����<�����~>ߏz���] -��*�U�<O�c2A��qX^�b��̭�����@DiwU�`�4K����;��;�=���XR8Vg"8\Hd|�RE&k�cOL�<fJ
�x��\n��3ŉ�us�Y\�Z��8G��i+K��Ҵipl��%i�O��y5�̐6is��b͔����C+�s�Z�]+"�Pa� �"f �Y�6�e��j)��?A� ��_�y�2����֯a�B"W��k�Cz*j�_��H�& $ϿEv!.��\^5!�*d��1�^���d!�Ǝ�D^�B<:,$\$"�U���<��ܚ���_9�o>���ٗ����jeK��,�4]�KH`&в皽�  w�J�vn[w�$�RrV�xTd<	����f׎�o��bU(
�`M
�U��D��d�
]�ɛ2�k�R8)_�����~�kK=F��7����Z9~2G�4�K�3*����������^����r|�grݸ���e�:�ʛv��#1�D���]���b��,�{_��D��� �����,���O&C[��ԃI��2�󭽸oIߏ�  1���T���������j.�F .�(F�+���>	�C���ū�{���&����Kp�%��������ut�.�	1��k @&�t����
-�C	h��D*�ٞMcge�Ir�f���%������m_�A5:��<zA�4˧�%�&�9p$��q2BRѪ�7I�B׸�$Xk���U��䊨)M�H���Lw;u�j�٩T����pLX ��`��i�m���� ���s	���>)��f�/Y���6�Bh����r0d�^P���xd����ӻN�����)d�+���و���M�H������a�z��5L����{p7X5dQV4��{�]�޶�w��)�s�<ׂo�{���إ����0"
�\��P�I������e^Ka�L��w�(W�	
���
����w��CG
"<R�JH$��D��]�Gw&���q7����G��s<1M�Ղ�>9����v�B����
��:Z[��'�iܒ��JYNiieR���  >��|U7Ԝ%��KN���T����@�]U!����"�bb����B���<8�� �?���tW	 �bY��R���K  R#+��L?@h �EV���28F��Ԧ�H �6L�P�i��p,X�Je!��r�h��վ��-��f��s�����}A
p�O�m�����]��]^n�IG~��u��\@��ݹ���"4
�-�@b�7)�ۧ���YU��=�� �
k�ݽ#�;ʷ�?j�9��*���=�\�NǠ��䜼e���55�"*U#��b��O��H��+�8.Q)e��R	� D$�%���M-����K�1zm��:3Ol��<�B��0B ��iMèi����-���+[��3��7��ׂ��AZ!��M �_���
0�p�gl0-�����I�˽w�|fR�->���;��O�;s��ݧ_������- ��0z.�t/�8�+�m�̙��h |@(,q�����#L�LBoH��
[N�L����v��^���G>4T7�	����[Ϟ�	����	$�������sBΪ��T*����dzIpx>.?�B�^��b	��;�v�F�;e��3�<�A��
��^���lT�<��xp�������r`da�,-_���m �o�l( ��x}�̒~*H���@ ���u��F_-{��&3�j9��������������������O�����/0%�s�X@<�)�/x0�=����צ0����- ) ���
`�G=�ܩ<Ɩx@�{�Ջ7�����z��� 09�0wp��M{|WNR5�J��H�p�x�Lr")')??W/�8^r�x��]��ʹ�l��5�hf�}Wf�:�>���d����Mz��U�QE���c#�  ����O�̼�)a����S�K����ߘ���N!<���
h�9�ˍu�K��JN� �H�
�:u�1����bEj*-99�Z��(-���FE]ͼ�y���'�1�&���w�W�r�
"�D"G���s�^����I�|�����!.8�����~�b�q��0�J$�HY��ݙ ]�3H�h�t�F�%��G�0�c��LNN���''�9�Q���E�rο&V��\釥9g߉���?�/�dTJ<�������9��C?�Y��s�S՚q`���E\��;��&�;������D'���t�Ts�RL)8$&D!?j�a&Q$ p�! ��@3$$!8�b�o�AI@��E\=���i��|�Dӹ���.y��.����������NH���-(�N�
kj&�� T���[,��á9(<�|��c=��*�:������%���E��˗ ��4!���*S&�q���:��#GNf��5;�رc���`���/�����?nOMM�l6|��nDv�ݔj���8 ��+@u�é�� ���ڧ�����Q�
����Փ1{�g�-C;�fK$�`�ݨxs*:
f�`�e������Ri�/*���{�R�C����T5pbERiEB@�ш����H��>�+(��o7*���i��>�L`��M��Q�!R5����>BT�d*{� ������O���e8G��~-^��g�u���ᚤ�@�_���I�����, �����  �L�4!�T*��C�1�Ri~���f��Ċn6����f��~�� >�����^����鈴}�����ɨ�3 n��3���tF���ᛙ[tt�r��$?`K)��đ(���;�%��kg$��D�G�;�H$
�!75qX��T�f���|�+>���"?�*>~ �������B>��mC'�Qv'j6(�	��/�7���ڦE ��w%an~����g�����&Sy�� ���_H��� u �zn���&���j�� < �O?v��%A+��    IDAT
�,�f�8��:�Aq�I\X(�D6�%�v��}X�}��O�zrÖ�U[6��G�ԣ,�|>Hc�%'
�X��|~!�2���k�T±{��I�.o��;����,q&֫=�<]}��*��b��H���'�3k3%A�,2�A�K,��E�dŃ([��4�t�T�֣9�_�G�J��&��އ|��lS������������ �w��18�)�D	4�Bw���:r,H���3�\�9�ۣ4�L � �=�������_|�<`�՚�z53:�X���p�)����fΒ�k�×ĝ�[�~�h+ 8�t~<��ޓ��U^�b�򬗞]��s�FT��=��v�}�o� y�/��	\�[�Kː�9�o۠NcQ���G	�e0:����=�Ÿo�Y^��+��S7n�����{�>��(�w�R:�#�TH�����֯[��'���8w�����k'Q�m'�Lβ{?xB"�X����!F�à3xl��4Q�u���Q�����`RR�-$ %@�?�(S������V=mBF׏�Pn٠�7�vG��A�0?oW�Y�7fT*Sh�|�,EU4��٧x���h�U���3�r2C;�8��<J�u�ј�/Hs 8�ǄJT���oC�*ڌm��(j�F�
9��ieoyoy9
� k�um�i���� ��#���]Y�:`d/�c�8����B�L��� @���cD{ũ���R�ޣ���n��y�� ƬX� J�vp8@��3Cl�*�[Ѕ�����/����U���X
d* �&q�|�*�A���R`����*��.�P���= ���.�;�P���i����r�`N��'�����>��n�V+b�
Űex~vnϞ=g�<����@�&:Z����F�"_8JeRɤ�X	c��R&��л*����<9]ƕG���[F��(akO2iC�O0���ЙP�0����N/7v��R#��@@��h1;���{݈^�|�����u�;a�r���:�k�f. �7�$ DR��%?Q
-�N�����֚�*�*��S��S��ߡCX����3����7*�+�ʌw2��ߠ,㻯��Q���s��gT�f�f�Գ�й�'J�H�4>�{������
�E[!#��������ՊN�� �vH[��XL2�-�H�}e�Q���#��&hhfr�酅��(���<�Á�����t*p�x��QȊyTj0�),�`�&�Ȗyn^���ps��~�w1�o�+ݽ|׹��\G�Wm^� �p�֏(N;�8�:)bC�؏��@��t��Aqwۧ1)��ŹG�F$�H���ई��1'L���#���թ�jQ��5U�w2o]�6��������
��&���
o�ba�Fi�U�]�!��ߣ[`)����[�d㿙���ZZZtvð�����՞�ϡ��D��ĵ��jA�����׍h�O���$����Z�Y� @��x��ba�&
xtm:�˅B��^����<��unބ�� �Eȥo��\���ܭ�:54�ժ��T*�Y �vT*����7w��0�s�H�K4��'l����}���-����:$+�m�	.�`�e�	� �E";�?��V0bG���\E�{�0G&�rsϝ+-�3�a���Tg|c��������_�P�OK��k:�\�,�G	��G�ݞx@7�w�_s�b�I�4.�V;�����[�súP�\�@���s���Y�SOý�	�! D���(,�Bz�Y�@�ىw@�TT���kK��|Ms_��Y�7��u�'&�����5yeq��e�X:ę�qT&�̰&3�"�L 6h� �A�#�B̀R�!nHp$%5M��:`�	��BQ*��JQ*.A���J���l���	Zwf?p�!O�o���9��{Ne�٠7��f=����;�/�,�������"*5	�"\.2� 
F B �O ��S�s���%J�p �=R���e�(�U}�|��S�z�oP�ȯ,�}>����E�p,"�eY)eَzMY�p%��4�F��)�e�����-�B~nn���s���&&��z��
&��d��@��wu������	~��	HT���H��_79L�s(7|K�jB�~x���?�{�7�%�� >�C �k��*��_��r����I^_��{���8t�NRh*�!�N���mci� {K`����M�X�rsA��hq�� ,�8�)5)I�����q�ZԜhcQ�N�H�0{�-��aa��d�!�b�^�?}��<HA�- '�@��4
�F�B��ʭ���__�M[#I[I�!xWRƙ�F���[	ޛ����Vg���~�ɧ[�E�������?0>0~�v��������n���qI�~ b��������<Jxt��-"ӏ3�d�ր�0���0&G�G�-�,?"�ea���`���@ �_�C�� ޳w'֜�rÜ�{��:G�V��j1�&��7U���?�G�8�M�� �,��
�Y��ݕ��I�틈8 �7�k�/RP�q =0rU@�� �O F�`*xY�V��<�O�	�v�#�f	����B�h�2�}���������E�V�k�ڵ��q�dj	G{���|*���MMv�����N;���k�����)���s�����G��X�@,�5�B�0-�'�(�p\��ha���8�Ņ�م�%@�8
9|�)!�`a�0��V^[�
���T>5��H��>�UM���V^^���:+<|����Q���┣��g*̌��a�a��I{�{}#z���9��<��#x��J�RnY�	��L��S!\�ⶱAL̠�M�AAH����S�?B@.�B����W�s |��"�"���Tη���{p�GB��8����ُ�?2m[�T79&i����	j/�?x4��������dQr˨�g�GD�]���e��Ǿ���+�
������gL7�u����yh1��LeueD�e���0�`bM�7��s�@��/�7_��Ĉཙ�|�����g��8��x�3�F�v�m.>��x� �
м���e
7�W����ş����G��o�xN�{&��Q#H]}1`;�!�����L� x�^ǅEt6��h�?ޗ�*l��JBBHX�8u!�s� �w6�$E
�z-۱�&  l4����n'>;v�S�$�������m���ퟷ�G��	[��5���^�Güp�y;��}�Ѱ��5G[a_���=�W����y[PJ�?�����]n4�!.��&�df� k��� ?`Yd%r�L>�q��@!X�4���t)JdLx���b 劒�������Dt:5���>i���S��]UVA4j�~3��Ù�)^�����K=]���Oe��^9�区YX�l��*��~�&�l	�Tg��&���a��`���5>>~�!����Y��X�� � �
�^�u.��d�)>	x#�����w�=���6�5�k�5�'n��>�y�f��l�x�QN�V{'���pNN�V[W]W��V��c���sk�sz�EsO����	��7��^~]�
���2dY�����BgE0�M#s�}@��e�1`RMTM�L'&/a�\�ӟ���QEcO����O��	VUi����B&Ia�$3%��K�T�ן��/t}sym	��vW����׾�Nq �.5Z����(tT)y�'A�=T7��|y������|_�8^��}��J��-�b�
�3 0��b^��pEG���A�:�v�'P
�D	P<
�BN��ђ��^���d�?�7�LK��3c�]�����#t�m�+5-�Ng$��5T*#�ud�j�m�ǡY���
ro� �� r����f چ�X@L/������A>S�|�bZ\pr:��� )�ʛ�L�q�l�A �6� !b�0ܘ���?S�����󆻇�yf��6�9�N�;p@�(�J��;{	C$�x[^�XϷ/ �>o����݊͂�ٚ�(S��/T9T}�!�5�5l�&eTd*I�C�� ��g�aI>��v�*�	��l׊����t�>66��T�	�|�F�!'!n�<�?�N
�4�L���յ$sӤ�1�1�6�	� ��oy�s�x����=-*zE9>|R/9x���ƨ(�c�t�C 1���`iR ���/�(��|F��X2�|~@Q.. �	�TX�H5��s��V��1X/&�T*�{�;���6vqK�:tTW�]p�P�n��*�(ظѫ!Z����O\���2h�D��X]Z�e$Dz
���½���4�R3����5��e�	��,s��#��{��oğ��!H(p-�,c ���L�H�: [�y�X6p�ظ�M��O���s�i:��8q���L��N�%�� �@�<+�I�6
�2���؂�(���K�|LK)T�-K�v@)�@)��@�V�<3HX&{�<
�+��$����m�?��sϽ�|O�G2��MHH@{x���R�/�A!���:�G��䋗�ɀ�dR/:$_>��x�4��|�)ᜇyV��@��A��Q�- ����C���H�˓������o��c5���9������H�8���i��wU@4�S�,8��8�����SI�ߊ�,'U
w�{
D,��f�$�6Cp�v�Dڥ[O�x�O&���s?�"\���L��A?��C̦�> �g+���kw�	d �ϸ�٩ ��_φ�&g�U]C��*}H��J�z��4���t��pD��b�GqN�[R�D�"�@n���Y����d,_B�p##����d"qr�"ʵ�x~8T__Zp0+_K=6��"�m���<�[��)dC>�d��b���3� E#^��A���#�2�P�a��f�8�o}��XZ��e�� �$Q���{�Z�W��Y�'�����V�m(+nx�iʾx�@�����I��~��e��,AѲH����a7���e{�[� ?{��o�]�v�N�tJѥ��w� ^Y�R��G��(ż��3�L��w�˳Q���U��Ƭ�_��]����ۓ����T�rn���H�B�/�w�6E���74��7���5���_����V�^.j��n���B{�t+C �[0�U�Jz�&yw���S2
 �e�0�Fp{���(ټ�t4��C7rxB�dJ�ogT�X����u�[---~1�����Ƣ����%�Rc��r�EE����R�D�pڢu+[���������[sj��×�+��
�)IԸ������p���T���_�5l�=���N�A�k[խ�?;'�X�`����w� ����PÚ�����u�����亠y\�!o?�����7$�f��Y�L�r�r��)E̓�h�ū�U%5RS�B+{PS��;��JL�݂�Ӄ����B���hz9�R��x�l q�d$�]l�/���h�`r�1��(�",�N��7{Ъ��HB����ꙥ_�}u޾8�����)(������I���48�<
�t�V�j�a2�#�=04m@�Ώ� ?�g��J���F��G�VRS�j�BjyyI,WB	���=N�H�pd��e[�{���4z���uԽ�� @F���<�� �K����5p�C�8�՝�ǹ�+}]SL<%��� e0��GKm#(��y����A��h7ML��ڧ�-���^�P�B��N�3��dj����Ů�'�^�v=�p���\Q���!�  �
� ���jG�Q"��� ��F�ca��F��%�M\mIʁݜ�p�̃��3�z G��>�gsZ�>��{2R�ר=@K�VJne���OO�nQ�����e~���bN�Ȫ�v�3�3�3g1�.&aO�9|�3��72(�bʻ�,���(��v�A����X��7���e}mui'h� t >4D����{��y�.�!�Q>v��Oie%���OT�耺�a���G=f5�*�d�����ۣ����L��t���EB"��1�T71!�I�q��o�R��C~xѕޒIZ|��B��vY�݌�jr�e V���$��|
�!�w3�Ř�VN�Ɏ�p�1�}��m0�; ,��Wݙ��k�{�����H�(�1 �lay�uV ����?�T�l�6py����퐫H�k"V�ȞD8����� $��		^��K̲e?��V��0������f�J ��q
����VV;�����,✦3#`�����a^��G������׈k�sZ�ʆ#�κLi��&�?�3Vs�% @:����]�Fu	�a(2X>&+R�njׇw��j�U>nx�Pp.[���?���%�ɼ��qf�Id�u^������k�YW���}��V�1/����.��z#�0���ā����ϝE��+�@�,^�0X���Tœ.�u�6<UwL�]�d� ���\^1�̅�xlQ��",:T�����Ve["���ݿV��Y�`P%���f��y���y�+����y�B��1�2�  �YėmF@��VI[V�Յ饬׊���FE�J�=6>�������2���r�������ƪ��Lw���d���s4�@�`�NW28�{�Vv)�2�t�dRo�B��|�a~yk̩fne�֣��Whi�k�����-��{�f�k���,��-�̬v� hp�bA�k���<�O8c���H����Z��ue���C ���2�<�t*���_PIˁ�~�. ��r�3����*D�6�k��k1(neV�&�������OcpN�!d^k<�r�� �Z���ԝ}Liǉn.'w*��aΗ��g�Q")^ڵ\l�]h�(�n${���������!�p��J9\�,��/hK�E�"ӡ��P�m���W%**�����=u�]�ä�癆@?�=���^�%��,�u\b4U'�Ȉכ��ۗ������].�F^�!&G��7/��n���gZ���vt�`�+s����k��I��P۩b�pP*�
�9!��寣�o��;!��zgg�`VRB��+.	W!�r�O�q�#��j@`�����Vo��F�]q����R����ǥ���y�O~U4�&d�wl�|�6�=S	�2���7�����>������EE]��`��)mWc|�j���u�&������Q[�y�5Z>�-'B뗜V\���!X��=m@[�L��e����)�mP�b-iu�C��Z6a���a�
��B1��32ʙVp=�����<5��>���R���g���A�������Tv�p	.#���+�� ���,l�6l����@Yx
���ŋEo�XM"Q'�5� diIq���`�JK��?p��I\�	޼�}�fޞ�{�ؔ}�?�3�V�Wۙ��2Y�hBx �h:u 
�J&��V� �`����7SS7oX^:a�s�ԕ��Z-�~>5f��?�!Ѡ��:�u�����
h���à���?����3�W��YY��+����N�qo�UN��3'�Ng��)٣��+{;{�>>������x�GTn�\���D0��u;~�g;y��M;�9��}�݆��_�?UII������24���W��@����E�돔��85���1�!9�;���L�RT~6�6�ߴ.�;���y�B������VVc�����
�I�O^�׳�վbi��ȱ����;��LO4�Y�:C�v�5����u��x��ȥ;J��%eO�4*@'˝t�/׆��;��!��&�d�FMM4����76�.T�I��l�:�j'�t�'D�_�O�U��9���,�D�m|�)`��X�[[�[C�E�|n�⺗��>]���"8��~8	��K�����hL�UЕ��eS���W���w�zy�֣	�Kw��{�
��Q��_��\���oh��cE�A�h���l�M��g��3 9�ņ�VL�-@\<L�#@X���>(�ŤA���u"��N$n8����r��<�:IL�p���3!6t��
p�W�Cp���ZP��_MF7�J�]�Xo�l
BI
��c���U���x�$�L�0�����h�5�4����L�E�v�؟$��k�Ū��x�  ���� B�[Q�N�9�h���g݆�E�U1��W�Hsv�D�\0R
Ʒ� �>�ЁN��I)��픆	�J$�[���&�PI��ߗd����$�\k�W5���O�=�%U�畯�ng�3{8��Jw{��9���E%��un��8��k�1U�n��`~���
�fPKF����ON���ʨ>_����ގ��q�{s���5D��'��~���Dg�28N���n�ҴY�K������F��S<����<�����?ςG�2�6R�[����f�~5�q��HF0���n˘>���J���q�Ͻ;����Gqt*Y/e�Y�t(U+A���/��,E~ˡ��X
0J+xN�F_�T4�PK�������S

0h5�X�($����7�:�C�t�5� �چ#���O��X1ykg���l�gMS�-�� �,�q��ӯa�P�6N�o>E9�6u:�(�B��0���������_�����d�4�U�OH��x��^$�^_��w�XǙ��N@��	j�8ҹ�[��i�t޾E}��_�$?��bE����M���5�א
H�}�j�}z2t�񠋆��L�"J�yn��I�����߹����7�o�B��-��<�_���WB$�Q�!�i$m��1%2#J�}��{I.�� ��u��*��
�P�SDj���.S�T��m�j��x9P}�!7��%}�u�)��J���?Zo$Y�D��hG' ��TV�A���M�އ\]�������oS'A���7{Ę�UP���v�^$�MT�v��H�#|cY'<آ���/L�}�E"�
��Qi)��Lܴ�2|��"%غ�����B��|�K��!���X�������3�^��6+oP�E����YE�:R�B�Xe-Ó�==��R򏝄z�-�-�	��e�N�, D ��_㘜<yF����[,|�Ǳ��KB����ȯ��k�4SJ%miK�缞�����a�Z��t�?ڶ6��?�p#m �@Y�������❶������V!�B�Î�m�4cz��p�̶�./�-���l���'F��ͅ{.�y���'���Ʊ�Ɗ#)��Ը5dez���K�"�gPy��[���k[ΠG�L�ZK���ѧ��'?a�_>|������9hDN�Ɖ%b(?�@�]˃�9�S�cI:���r�'l���}��~ۍ�e������z1)s+t|7��k��t?�еʹ��ؙ5p��i�d�a�t���,�GJj��*߯_�%�F�ξk~�sշ����n�B�����X�'>����f%�U�~7o1��?�@�?�7���"朗��؃���	�>��w]-T�iɵz�q@�2ZXr��@j�������̹r4/w��-[<�a$�Ul�]��m��;��%IC2c6��K�]���:����&\��qdO�K��[�Οa�)ZK������<ou��֖Zڵ蠛K���9���l��bneCU@�	>�,�x�8�`n����/��� �#�x�9��o^��0Oys�N�﹑~||<ֻ0�/�����ۼ�lu��X�����$�C�R�1��O�W��9�8���A��Z�7~���qk�t���'�\|WKK�c�/��qһju�=!]�Q��|-3�2����ڪ�38�
%��{����%$���ɣ�x�@�x8�Ơ8<�;����ǉ����g�_F�
**��� u�q��TG~m��1F��W�4myz�S���B�_�o6uG�����~���Z^c�&ūm��� �1���/m�"cZۋiڒL��B�·e��p�%~���41-냯W����]�`�bR���EX)�z���t�2��I3������s�⋎�[k����{�v�:(�!:d�����u	���������lN��-����n'��@;���`�f���}=�_<���W*<�����
��>��)灚�����d]aL�;y�]L�7\g�6'�S1,��Bl��P=}�QD1�ژ�]NP�፳�]2�����^��'P���㙴�ލ{$�HG�0*"^?"���r�]q��qἕ{��
b����52<N8�wų$;@@!�7ٵ~sk�{2�KF�>/�F6��wv&]d��ID��rW�_�^c�lQ?�l2��Ę=�d^.�\)b�肹���y>��ΛN�25�=�MR��ߝ(Sq��o4�>�|���ö� �DL�?=�KJ`P��l01P�8dN���������ڦ��k��i����m�|�G�a&R����47Wg�hlq��M:�Dա��bad�*�J~�f���z�7bҫ$��s���}1�ur�?�wu�UR�Dڜ���/p���F�)�,s����sT(6���;�bske��)�pe�u�O��$��ʈ��;J�$��R��6��#飃_��WT�K������5��w��#���&�m�7A�����¬Iص,�k�3����O��j���,�'C:3o��	.�~)}uq�t�ٷO�Oֿ��N��f[������f�+7�i�.7����-�>��Z�*�C`�m��;7�"�`�j��fR�4x2m�`�4Ӓ��<��n�	����|���4n�_2�l��{���_�T�Gf����%^v!2ɘ-e/��b���w�������x�~��=81�5��ndP����m���f���`�]�p�WgZH�\��}s�Q��H\Z�bK/_6��4��Uw�K�2G�n�|��C.[~��f������R��6�ݙ�1�j�۾����=�:���U/i}cҐ%����ΰ��</�����7�ul9%d|���6Ȱ���w\1�~��1u�`�3X5������`Eֿ����Q�
�O�O#,[�$��Ln$��ޒ�Ӝ]?�u�$�6��5���	�d���%�*q��6%�<a����׽�<��=�y�`��}���o6��Ԯĥs0�{!Í2��Z�ey@Ou����rpU�l�Y�Sg;h���!�
��p�t�uӌ8Vy�Qu��[�o3~
�!��qSE�/j�s�T��;�v�r�R�9����a�����VrITB3o���ԍ�cW��;�)�ח�����Ӓo��n���b�kҋ>QZ�ң,�h^I�mݍڒ�U�C�ss_r�L0���$V��u$o"���p��f��]^�,����-�z .~v|�M�"���+����ǰ�`�¦(�����5벌��baA4|�袰�-����Ί7�
�q��u��J~��)��a^S�\w�b�����ښ�4J�߄�PK   ��W��2�o       jsons/user_defined.json��j�0�_%�lI�זo����R�s*�8��
ɕ���]'Mq���&ig?�.�%ݦU$'�W�R�6�"yW�kk��(�_|��������X�3S�©j���M�C}Ytji���	��'|]aWi��L�4��a!k�:ͤ*��3;���՗����mw��m�N�g�ik���j�#X�o��WS�ۦ�\�g%<��2�(�����I���F��h�̪��i��
��zpz�|I$e��<H�QH�=C�+S�Z���I�b�=�?���J� ��"�O�u��s�b��)�h�A!$�ȑ�s���:��g"
�eq
�����?2��B���ζ�uz��!o�5L�����K��y��PK   ��W�� ��0  ��            ��    cirkitFile.jsonPK   ��W`�����  (�  /           ��1  images/a675022d-8297-46f2-a9f0-ef789ec00656.pngPK   ��W��2�o               ��/ jsons/user_defined.jsonPK      �   �   